-- megafunction wizard: %ALTASMI_PARALLEL%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: ALTASMI_PARALLEL 

-- ============================================================
-- File Name: asmicont.vhd
-- Megafunction Name(s):
-- 			ALTASMI_PARALLEL
--
-- Simulation Library Files(s):
-- 			
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 18.1.0 Build 625 09/12/2018 SJ Lite Edition
-- ************************************************************


--Copyright (C) 2018  Intel Corporation. All rights reserved.
--Your use of Intel Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Intel Program License 
--Subscription Agreement, the Intel Quartus Prime License Agreement,
--the Intel FPGA IP License Agreement, or other applicable license
--agreement, including, without limitation, that your use is for
--the sole purpose of programming logic devices manufactured by
--Intel and sold by Intel or its authorized distributors.  Please
--refer to the applicable agreement for further details.


--altasmi_parallel CBX_AUTO_BLACKBOX="ALL" DATA_WIDTH="STANDARD" DEVICE_FAMILY="Cyclone V" ENABLE_SIM="FALSE" EPCS_TYPE="EPCS64" FLASH_RSTPIN="FALSE" PAGE_SIZE=1 PORT_BULK_ERASE="PORT_UNUSED" PORT_DIE_ERASE="PORT_UNUSED" PORT_EN4B_ADDR="PORT_UNUSED" PORT_EX4B_ADDR="PORT_UNUSED" PORT_FAST_READ="PORT_UNUSED" PORT_ILLEGAL_ERASE="PORT_UNUSED" PORT_ILLEGAL_WRITE="PORT_UNUSED" PORT_RDID_OUT="PORT_UNUSED" PORT_READ_ADDRESS="PORT_USED" PORT_READ_DUMMYCLK="PORT_UNUSED" PORT_READ_RDID="PORT_UNUSED" PORT_READ_SID="PORT_UNUSED" PORT_READ_STATUS="PORT_UNUSED" PORT_SECTOR_ERASE="PORT_UNUSED" PORT_SECTOR_PROTECT="PORT_UNUSED" PORT_SHIFT_BYTES="PORT_UNUSED" PORT_WREN="PORT_UNUSED" PORT_WRITE="PORT_UNUSED" USE_ASMIBLOCK="ON" USE_EAB="ON" WRITE_DUMMY_CLK=0 addr busy clkin data_valid dataout rden read read_address reset INTENDED_DEVICE_FAMILY="Cyclone V" ALTERA_INTERNAL_OPTIONS=SUPPRESS_DA_RULE_INTERNAL=C106
--VERSION_BEGIN 18.1 cbx_a_gray2bin 2018:09:12:13:04:24:SJ cbx_a_graycounter 2018:09:12:13:04:24:SJ cbx_altasmi_parallel 2018:09:12:13:04:24:SJ cbx_altdpram 2018:09:12:13:04:24:SJ cbx_altera_counter 2018:09:12:13:04:24:SJ cbx_altera_syncram 2018:09:12:13:04:24:SJ cbx_altera_syncram_nd_impl 2018:09:12:13:04:24:SJ cbx_altsyncram 2018:09:12:13:04:24:SJ cbx_arriav 2018:09:12:13:04:23:SJ cbx_cyclone 2018:09:12:13:04:24:SJ cbx_cycloneii 2018:09:12:13:04:24:SJ cbx_fifo_common 2018:09:12:13:04:24:SJ cbx_lpm_add_sub 2018:09:12:13:04:24:SJ cbx_lpm_compare 2018:09:12:13:04:24:SJ cbx_lpm_counter 2018:09:12:13:04:24:SJ cbx_lpm_decode 2018:09:12:13:04:24:SJ cbx_lpm_mux 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ cbx_nadder 2018:09:12:13:04:24:SJ cbx_nightfury 2018:09:12:13:04:24:SJ cbx_scfifo 2018:09:12:13:04:24:SJ cbx_stratix 2018:09:12:13:04:24:SJ cbx_stratixii 2018:09:12:13:04:24:SJ cbx_stratixiii 2018:09:12:13:04:24:SJ cbx_stratixv 2018:09:12:13:04:24:SJ cbx_util_mgl 2018:09:12:13:04:24:SJ cbx_zippleback 2018:09:12:13:04:24:SJ  VERSION_END

 LIBRARY altera_mf;
 USE altera_mf.all;

 LIBRARY cyclonev;
 USE cyclonev.all;

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = a_graycounter 3 cyclonev_asmiblock 1 lpm_counter 1 lut 6 mux21 1 reg 91 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  asmicont_altasmi_parallel_ehl2 IS 
	 PORT 
	 ( 
		 addr	:	IN  STD_LOGIC_VECTOR (23 DOWNTO 0);
		 busy	:	OUT  STD_LOGIC;
		 clkin	:	IN  STD_LOGIC;
		 data_valid	:	OUT  STD_LOGIC;
		 dataout	:	OUT  STD_LOGIC_VECTOR (7 DOWNTO 0);
		 rden	:	IN  STD_LOGIC;
		 read	:	IN  STD_LOGIC := '0';
		 read_address	:	OUT  STD_LOGIC_VECTOR (23 DOWNTO 0);
		 reset	:	IN  STD_LOGIC := '0'
	 ); 
 END asmicont_altasmi_parallel_ehl2;

 ARCHITECTURE RTL OF asmicont_altasmi_parallel_ehl2 IS

	 ATTRIBUTE synthesis_clearbox : natural;
	 ATTRIBUTE synthesis_clearbox OF RTL : ARCHITECTURE IS 2;
	 ATTRIBUTE ALTERA_ATTRIBUTE : string;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF RTL : ARCHITECTURE IS "SUPPRESS_DA_RULE_INTERNAL=C106";

	 SIGNAL  wire_addbyte_cntr_w_lg_w_q_range140w145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addbyte_cntr_w_lg_w_q_range143w144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addbyte_cntr_clk_en	:	STD_LOGIC;
	 SIGNAL  wire_stage_cntr_w139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addbyte_cntr_clock	:	STD_LOGIC;
	 SIGNAL  wire_addbyte_cntr_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_addbyte_cntr_sclr	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_end_operation90w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addbyte_cntr_w_q_range143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addbyte_cntr_w_q_range140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_gen_cntr_w_lg_w_q_range103w104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_gen_cntr_w_lg_w_q_range101w102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_gen_cntr_clk_en	:	STD_LOGIC;
	 SIGNAL  wire_w32w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_gen_cntr_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_gen_cntr_sclr	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_end1_cyc_reg_in_wire33w34w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_gen_cntr_w_q_range101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_gen_cntr_w_q_range103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w342w343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w342w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w347w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range93w96w339w340w341w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range93w96w344w345w346w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range93w94w95w353w354w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range93w98w429w430w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range93w96w339w340w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range93w96w364w365w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range93w96w344w345w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range93w94w95w353w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range93w98w429w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range93w96w339w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range93w96w364w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range93w96w344w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range93w96w136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range93w96w337w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range92w97w115w116w117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range92w97w115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range93w94w95w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_q_range93w98w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_q_range93w96w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range92w97w115w116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_q_range92w97w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_q_range93w94w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_clk_en	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_w_lg_w86w87w88w89w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_sclr	:	STD_LOGIC;
	 SIGNAL  wire_stage_cntr_w_q_range92w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_q_range93w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_sd2_data1in	:	STD_LOGIC;
	 SIGNAL  wire_vcc	:	STD_LOGIC;
	 SIGNAL	 add_msb_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_add_msb_reg_ena	:	STD_LOGIC;
	 SIGNAL	 add_rollover_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_addr_reg_d	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL	 addr_reg	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_addr_reg_ena	:	STD_LOGIC_VECTOR(23 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_q_range403w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL	 wire_asmi_opcode_reg_d	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL	 asmi_opcode_reg	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_asmi_opcode_reg_ena	:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	 SIGNAL  wire_asmi_opcode_reg_w_q_range150w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL	 busy_det_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 clr_read_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 clr_read_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dvalid_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_dvalid_reg_ena	:	STD_LOGIC;
	 SIGNAL	 wire_dvalid_reg_sclr	:	STD_LOGIC;
	 SIGNAL	 dvalid_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 end1_cyc_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 end1_cyc_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 end_op_hdlyreg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 end_op_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 end_rbyte_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_end_rbyte_reg_ena	:	STD_LOGIC;
	 SIGNAL	 wire_end_rbyte_reg_sclr	:	STD_LOGIC;
	 SIGNAL	 end_read_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 ncs_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_ncs_reg_sclr	:	STD_LOGIC;
	 SIGNAL  wire_ncs_reg_w_lg_q390w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 wire_read_add_reg_d	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL	 read_add_reg	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_read_add_reg_ena	:	STD_LOGIC_VECTOR(23 DOWNTO 0);
	 SIGNAL	 wire_read_data_reg_d	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL	 read_data_reg	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_read_data_reg_ena	:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	 SIGNAL	 wire_read_dout_reg_d	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL	 read_dout_reg	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_read_dout_reg_ena	:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	 SIGNAL	 read_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_read_reg_ena	:	STD_LOGIC;
	 SIGNAL	 shift_op_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 stage2_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 stage3_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 stage4_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_read_add_cntr_clk_en	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_w_lg_rden_wire491w492w493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_read_add_cntr_data	:	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  wire_read_add_cntr_q	:	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  wire_read_add_cntr_sload	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_rden_wire491w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	wire_mux211_dataout	:	STD_LOGIC;
	 SIGNAL  wire_w269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w209w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w202w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w485w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode166w167w168w253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode166w167w168w169w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode171w172w173w255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode171w172w173w174w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode205w206w207w208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode176w177w178w257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode176w177w178w179w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode217w218w219w275w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode217w218w219w220w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode198w199w200w201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_read369w370w371w372w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_read301w482w483w484w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_sec_erase44w425w426w427w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode166w167w168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode171w172w173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode181w186w261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode181w186w187w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode181w182w259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode181w182w183w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode205w206w207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode176w177w178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode217w218w219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode198w199w200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_read369w370w371w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_read369w370w428w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_read301w482w483w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_sec_erase44w425w426w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_4baddr158w159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_ex4baddr153w154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_write189w190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_write53w348w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_end_read_byte489w501w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode160w249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode160w161w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode155w247w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode155w156w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode191w263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode191w192w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode166w167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode171w172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode211w271w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode211w212w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode214w273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode214w215w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode194w265w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode194w195w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode222w277w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode222w223w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode225w279w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode225w226w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode181w186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode181w182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode205w206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode176w177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode217w218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode163w251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode163w164w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode198w199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_stage3_wire35w36w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_start_poll355w356w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read369w370w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_write62w110w111w112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_write62w63w417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read301w482w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_sec_erase44w425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_rden_wire421w422w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_addr_overdie412w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_addr_overdie402w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_4baddr158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_bulk_erase349w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_ex4baddr153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read_nonvolatile335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_write189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_write60w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_write53w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_operation520w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_read_byte489w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_in_operation28w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_not_busy414w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_not_busy406w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_opcode151w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage3_wire419w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage3_wire311w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage3_wire449w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage3_wire300w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage3_wire45w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage3_wire35w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage3_wire404w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage4_wire451w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage4_wire302w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage4_wire420w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage4_wire316w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_start_poll355w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_write53w367w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_stage4_wire316w317w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_stage4_wire302w303w304w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_read_stat312w313w314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_addr_overdie514w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_busy_wire1w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_clkin_wire91w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_clr_rstat_wire26w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_clr_sid_wire25w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_fast_read368w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_memadd434w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_polling185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read369w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read_rdid41w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read_stat42w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read_volatile197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_wren43w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_write_volatile204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_add_cycle73w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_fast_read67w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_operation500w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_ophdly27w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_pgwr_data52w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_read70w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rden_wire516w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_rdid_wire7w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_sid_wire6w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_sec_protect_wire5w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_st_busy_wire107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_pagewr_buf_not_empty_range58w59w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode225w279w280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode225w226w227w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_write62w63w417w418w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_rden_wire421w422w423w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_not_busy414w415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_not_busy406w407w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_stage4_wire451w452w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_stage4_wire302w303w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode225w279w280w281w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode225w226w227w228w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_rden_wire421w422w423w424w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_not_busy406w407w408w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w282w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w229w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w282w283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w229w230w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w282w283w284w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w229w230w231w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w282w283w284w285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w229w230w231w232w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w282w283w284w285w286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w229w230w231w232w233w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w282w283w284w285w286w287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w229w230w231w232w233w234w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w288w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w235w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w288w289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w235w236w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w288w289w290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w235w236w237w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w288w289w290w291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w235w236w237w238w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w288w289w290w291w292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w235w236w237w238w239w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w288w289w290w291w292w293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w235w236w237w238w239w240w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w294w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w241w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w294w295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w241w242w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w241w242w243w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w133w134w135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w133w134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_read301w437w438w439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_read_sid129w130w131w132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_read301w437w438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_read_sid129w130w131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_read_stat308w309w310w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_read_stat308w447w448w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_write62w110w111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read301w450w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read301w437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read_rdid298w299w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read_sid129w130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read_stat312w313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read_stat308w309w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read_stat308w447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_write62w110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_write62w63w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_data0out_wire454w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_4baddr351w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_ex4baddr350w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read_rdid298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read_sid129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read_stat312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read_stat305w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read_stat308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_sec_erase44w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_wren352w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_write62w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rden_wire421w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  add_rollover :	STD_LOGIC;
	 SIGNAL  addr_overdie :	STD_LOGIC;
	 SIGNAL  addr_overdie_pos :	STD_LOGIC;
	 SIGNAL  addr_reg_overdie :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  b4addr_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  berase_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  busy_wire :	STD_LOGIC;
	 SIGNAL  clkin_wire :	STD_LOGIC;
	 SIGNAL  clr_addmsb_wire :	STD_LOGIC;
	 SIGNAL  clr_endrbyte_wire :	STD_LOGIC;
	 SIGNAL  clr_read_wire :	STD_LOGIC;
	 SIGNAL  clr_read_wire2 :	STD_LOGIC;
	 SIGNAL  clr_rstat_wire :	STD_LOGIC;
	 SIGNAL  clr_sid_wire :	STD_LOGIC;
	 SIGNAL  clr_write_wire2 :	STD_LOGIC;
	 SIGNAL  data0out_wire :	STD_LOGIC;
	 SIGNAL  data_valid_wire :	STD_LOGIC;
	 SIGNAL  dataoe_wire :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  dataout_wire :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  derase_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  do_4baddr :	STD_LOGIC;
	 SIGNAL  do_bulk_erase :	STD_LOGIC;
	 SIGNAL  do_die_erase :	STD_LOGIC;
	 SIGNAL  do_ex4baddr :	STD_LOGIC;
	 SIGNAL  do_fast_read :	STD_LOGIC;
	 SIGNAL  do_fread_epcq :	STD_LOGIC;
	 SIGNAL  do_freadwrv_polling :	STD_LOGIC;
	 SIGNAL  do_memadd :	STD_LOGIC;
	 SIGNAL  do_polling :	STD_LOGIC;
	 SIGNAL  do_read :	STD_LOGIC;
	 SIGNAL  do_read_nonvolatile :	STD_LOGIC;
	 SIGNAL  do_read_rdid :	STD_LOGIC;
	 SIGNAL  do_read_sid :	STD_LOGIC;
	 SIGNAL  do_read_stat :	STD_LOGIC;
	 SIGNAL  do_read_volatile :	STD_LOGIC;
	 SIGNAL  do_sec_erase :	STD_LOGIC;
	 SIGNAL  do_sec_prot :	STD_LOGIC;
	 SIGNAL  do_sprot_polling :	STD_LOGIC;
	 SIGNAL  do_wait_dummyclk :	STD_LOGIC;
	 SIGNAL  do_wren :	STD_LOGIC;
	 SIGNAL  do_write :	STD_LOGIC;
	 SIGNAL  do_write_polling :	STD_LOGIC;
	 SIGNAL  do_write_volatile :	STD_LOGIC;
	 SIGNAL  end1_cyc_gen_cntr_wire :	STD_LOGIC;
	 SIGNAL  end1_cyc_normal_in_wire :	STD_LOGIC;
	 SIGNAL  end1_cyc_reg_in_wire :	STD_LOGIC;
	 SIGNAL  end_add_cycle :	STD_LOGIC;
	 SIGNAL  end_add_cycle_mux_datab_wire :	STD_LOGIC;
	 SIGNAL  end_fast_read :	STD_LOGIC;
	 SIGNAL  end_one_cyc_pos :	STD_LOGIC;
	 SIGNAL  end_one_cycle :	STD_LOGIC;
	 SIGNAL  end_op_wire :	STD_LOGIC;
	 SIGNAL  end_operation :	STD_LOGIC;
	 SIGNAL  end_ophdly :	STD_LOGIC;
	 SIGNAL  end_pgwr_data :	STD_LOGIC;
	 SIGNAL  end_read :	STD_LOGIC;
	 SIGNAL  end_read_byte :	STD_LOGIC;
	 SIGNAL  exb4addr_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  fast_read_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  freadwrv_sdoin :	STD_LOGIC;
	 SIGNAL  in_operation :	STD_LOGIC;
	 SIGNAL  load_opcode :	STD_LOGIC;
	 SIGNAL  memadd_sdoin :	STD_LOGIC;
	 SIGNAL  ncs_reg_ena_wire :	STD_LOGIC;
	 SIGNAL  not_busy :	STD_LOGIC;
	 SIGNAL  oe_wire :	STD_LOGIC;
	 SIGNAL  pagewr_buf_not_empty :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  rden_wire :	STD_LOGIC;
	 SIGNAL  rdid_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  rdummyclk_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  read_data_reg_in_wire :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  read_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  read_rdid_wire :	STD_LOGIC;
	 SIGNAL  read_sid_wire :	STD_LOGIC;
	 SIGNAL  read_wire :	STD_LOGIC;
	 SIGNAL  rflagstat_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  rnvdummyclk_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  rsid_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  rsid_sdoin :	STD_LOGIC;
	 SIGNAL  rstat_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  scein_wire :	STD_LOGIC;
	 SIGNAL  sdoin_wire :	STD_LOGIC;
	 SIGNAL  sec_protect_wire :	STD_LOGIC;
	 SIGNAL  secprot_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  secprot_sdoin :	STD_LOGIC;
	 SIGNAL  serase_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  shift_opcode :	STD_LOGIC;
	 SIGNAL  shift_opdata :	STD_LOGIC;
	 SIGNAL  shift_pgwr_data :	STD_LOGIC;
	 SIGNAL  st_busy_wire :	STD_LOGIC;
	 SIGNAL  stage2_wire :	STD_LOGIC;
	 SIGNAL  stage3_wire :	STD_LOGIC;
	 SIGNAL  stage4_wire :	STD_LOGIC;
	 SIGNAL  start_frpoll :	STD_LOGIC;
	 SIGNAL  start_poll :	STD_LOGIC;
	 SIGNAL  start_sppoll :	STD_LOGIC;
	 SIGNAL  start_wrpoll :	STD_LOGIC;
	 SIGNAL  to_sdoin_wire :	STD_LOGIC;
	 SIGNAL  wren_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wren_wire :	STD_LOGIC;
	 SIGNAL  write_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  write_prot_true :	STD_LOGIC;
	 SIGNAL  write_sdoin :	STD_LOGIC;
	 SIGNAL  wrvolatile_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_addr_range413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_addr_range405w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_addr_reg_overdie_range411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_addr_reg_overdie_range401w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_b4addr_opcode_range248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_b4addr_opcode_range157w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_berase_opcode_range252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_berase_opcode_range165w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_dataout_wire_range453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_derase_opcode_range254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_derase_opcode_range170w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_exb4addr_opcode_range246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exb4addr_opcode_range152w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_fast_read_opcode_range270w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_fast_read_opcode_range210w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_pagewr_buf_not_empty_range58w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rdid_opcode_range276w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rdid_opcode_range221w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_rdummyclk_opcode_range268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rdummyclk_opcode_range203w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_read_opcode_range272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_read_opcode_range213w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_rflagstat_opcode_range258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rflagstat_opcode_range180w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_rnvdummyclk_opcode_range264w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rnvdummyclk_opcode_range193w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_rsid_opcode_range278w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rsid_opcode_range224w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_rstat_opcode_range260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rstat_opcode_range184w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_secprot_opcode_range274w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_secprot_opcode_range216w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_serase_opcode_range256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_serase_opcode_range175w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_wren_opcode_range250w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_wren_opcode_range162w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_write_opcode_range262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_write_opcode_range188w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_wrvolatile_opcode_range266w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_wrvolatile_opcode_range196w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 COMPONENT  a_graycounter
	 GENERIC 
	 (
		PVALUE	:	NATURAL := 0;
		WIDTH	:	NATURAL := 8;
		lpm_type	:	STRING := "a_graycounter"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clk_en	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC;
		cnt_en	:	IN STD_LOGIC := '1';
		q	:	OUT STD_LOGIC_VECTOR(width-1 DOWNTO 0);
		qbin	:	OUT STD_LOGIC_VECTOR(width-1 DOWNTO 0);
		sclr	:	IN STD_LOGIC := '0';
		updown	:	IN STD_LOGIC := '1'
	 ); 
	 END COMPONENT;
	 COMPONENT  cyclonev_asmiblock
	 GENERIC 
	 (
		enable_sim	:	STRING := "false";
		lpm_type	:	STRING := "cyclonev_asmiblock"
	 );
	 PORT
	 ( 
		data0in	:	OUT STD_LOGIC;
		data0oe	:	IN STD_LOGIC := '0';
		data0out	:	IN STD_LOGIC := '0';
		data1in	:	OUT STD_LOGIC;
		data1oe	:	IN STD_LOGIC := '0';
		data1out	:	IN STD_LOGIC := '0';
		data2in	:	OUT STD_LOGIC;
		data2oe	:	IN STD_LOGIC := '0';
		data2out	:	IN STD_LOGIC := '0';
		data3in	:	OUT STD_LOGIC;
		data3oe	:	IN STD_LOGIC := '0';
		data3out	:	IN STD_LOGIC := '0';
		dclk	:	IN STD_LOGIC := '0';
		oe	:	IN STD_LOGIC := '0';
		sce	:	IN STD_LOGIC := '0';
		spidatain	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		spidataout	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		spidclk	:	OUT STD_LOGIC;
		spisce	:	OUT STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_counter
	 GENERIC 
	 (
		lpm_avalue	:	STRING := "0";
		lpm_direction	:	STRING := "DEFAULT";
		lpm_modulus	:	NATURAL := 0;
		lpm_port_updown	:	STRING := "PORT_CONNECTIVITY";
		lpm_pvalue	:	STRING := "0";
		lpm_svalue	:	STRING := "0";
		lpm_width	:	NATURAL;
		lpm_type	:	STRING := "lpm_counter"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aload	:	IN STD_LOGIC := '0';
		aset	:	IN STD_LOGIC := '0';
		cin	:	IN STD_LOGIC := '1';
		clk_en	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC;
		cnt_en	:	IN STD_LOGIC := '1';
		cout	:	OUT STD_LOGIC;
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		eq	:	OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		sclr	:	IN STD_LOGIC := '0';
		sload	:	IN STD_LOGIC := '0';
		sset	:	IN STD_LOGIC := '0';
		updown	:	IN STD_LOGIC := '1'
	 ); 
	 END COMPONENT;
 BEGIN

	wire_vcc <= '1';
	wire_w269w(0) <= wire_w_lg_w_lg_w_lg_w_lg_load_opcode205w206w207w208w(0) AND wire_w_rdummyclk_opcode_range268w(0);
	loop0 : FOR i IN 0 TO 6 GENERATE 
		wire_w209w(i) <= wire_w_lg_w_lg_w_lg_w_lg_load_opcode205w206w207w208w(0) AND wire_w_rdummyclk_opcode_range203w(i);
	END GENERATE loop0;
	wire_w267w(0) <= wire_w_lg_w_lg_w_lg_w_lg_load_opcode198w199w200w201w(0) AND wire_w_wrvolatile_opcode_range266w(0);
	loop1 : FOR i IN 0 TO 6 GENERATE 
		wire_w202w(i) <= wire_w_lg_w_lg_w_lg_w_lg_load_opcode198w199w200w201w(0) AND wire_w_wrvolatile_opcode_range196w(i);
	END GENERATE loop1;
	wire_w485w(0) <= wire_w_lg_w_lg_w_lg_w_lg_do_read301w482w483w484w(0) AND end_read_byte;
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode166w167w168w253w(0) <= wire_w_lg_w_lg_w_lg_load_opcode166w167w168w(0) AND wire_w_berase_opcode_range252w(0);
	loop2 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_load_opcode166w167w168w169w(i) <= wire_w_lg_w_lg_w_lg_load_opcode166w167w168w(0) AND wire_w_berase_opcode_range165w(i);
	END GENERATE loop2;
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode171w172w173w255w(0) <= wire_w_lg_w_lg_w_lg_load_opcode171w172w173w(0) AND wire_w_derase_opcode_range254w(0);
	loop3 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_load_opcode171w172w173w174w(i) <= wire_w_lg_w_lg_w_lg_load_opcode171w172w173w(0) AND wire_w_derase_opcode_range170w(i);
	END GENERATE loop3;
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode205w206w207w208w(0) <= wire_w_lg_w_lg_w_lg_load_opcode205w206w207w(0) AND wire_w_lg_do_read_stat42w(0);
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode176w177w178w257w(0) <= wire_w_lg_w_lg_w_lg_load_opcode176w177w178w(0) AND wire_w_serase_opcode_range256w(0);
	loop4 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_load_opcode176w177w178w179w(i) <= wire_w_lg_w_lg_w_lg_load_opcode176w177w178w(0) AND wire_w_serase_opcode_range175w(i);
	END GENERATE loop4;
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode217w218w219w275w(0) <= wire_w_lg_w_lg_w_lg_load_opcode217w218w219w(0) AND wire_w_secprot_opcode_range274w(0);
	loop5 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_load_opcode217w218w219w220w(i) <= wire_w_lg_w_lg_w_lg_load_opcode217w218w219w(0) AND wire_w_secprot_opcode_range216w(i);
	END GENERATE loop5;
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode198w199w200w201w(0) <= wire_w_lg_w_lg_w_lg_load_opcode198w199w200w(0) AND wire_w_lg_do_read_stat42w(0);
	wire_w_lg_w_lg_w_lg_w_lg_do_read369w370w371w372w(0) <= wire_w_lg_w_lg_w_lg_do_read369w370w371w(0) AND end_one_cycle;
	wire_w_lg_w_lg_w_lg_w_lg_do_read301w482w483w484w(0) <= wire_w_lg_w_lg_w_lg_do_read301w482w483w(0) AND end_one_cyc_pos;
	wire_w_lg_w_lg_w_lg_w_lg_do_sec_erase44w425w426w427w(0) <= wire_w_lg_w_lg_w_lg_do_sec_erase44w425w426w(0) AND end_operation;
	wire_w_lg_w_lg_w_lg_load_opcode166w167w168w(0) <= wire_w_lg_w_lg_load_opcode166w167w(0) AND wire_w_lg_do_read_stat42w(0);
	wire_w_lg_w_lg_w_lg_load_opcode171w172w173w(0) <= wire_w_lg_w_lg_load_opcode171w172w(0) AND wire_w_lg_do_read_stat42w(0);
	wire_w_lg_w_lg_w_lg_load_opcode181w186w261w(0) <= wire_w_lg_w_lg_load_opcode181w186w(0) AND wire_w_rstat_opcode_range260w(0);
	loop6 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_load_opcode181w186w187w(i) <= wire_w_lg_w_lg_load_opcode181w186w(0) AND wire_w_rstat_opcode_range184w(i);
	END GENERATE loop6;
	wire_w_lg_w_lg_w_lg_load_opcode181w182w259w(0) <= wire_w_lg_w_lg_load_opcode181w182w(0) AND wire_w_rflagstat_opcode_range258w(0);
	loop7 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_load_opcode181w182w183w(i) <= wire_w_lg_w_lg_load_opcode181w182w(0) AND wire_w_rflagstat_opcode_range180w(i);
	END GENERATE loop7;
	wire_w_lg_w_lg_w_lg_load_opcode205w206w207w(0) <= wire_w_lg_w_lg_load_opcode205w206w(0) AND wire_w_lg_do_wren43w(0);
	wire_w_lg_w_lg_w_lg_load_opcode176w177w178w(0) <= wire_w_lg_w_lg_load_opcode176w177w(0) AND wire_w_lg_do_read_stat42w(0);
	wire_w_lg_w_lg_w_lg_load_opcode217w218w219w(0) <= wire_w_lg_w_lg_load_opcode217w218w(0) AND wire_w_lg_do_read_stat42w(0);
	wire_w_lg_w_lg_w_lg_load_opcode198w199w200w(0) <= wire_w_lg_w_lg_load_opcode198w199w(0) AND wire_w_lg_do_wren43w(0);
	wire_w_lg_w_lg_w_lg_do_read369w370w371w(0) <= wire_w_lg_w_lg_do_read369w370w(0) AND wire_w_lg_w_lg_do_write53w367w(0);
	wire_w_lg_w_lg_w_lg_do_read369w370w428w(0) <= wire_w_lg_w_lg_do_read369w370w(0) AND clr_write_wire2;
	wire_w_lg_w_lg_w_lg_do_read301w482w483w(0) <= wire_w_lg_w_lg_do_read301w482w(0) AND wire_stage_cntr_w_lg_w_q_range92w97w(0);
	wire_w_lg_w_lg_w_lg_do_sec_erase44w425w426w(0) <= wire_w_lg_w_lg_do_sec_erase44w425w(0) AND wire_w_lg_do_read_stat42w(0);
	wire_w_lg_w_lg_do_4baddr158w159w(0) <= wire_w_lg_do_4baddr158w(0) AND wire_w_lg_do_wren43w(0);
	wire_w_lg_w_lg_do_ex4baddr153w154w(0) <= wire_w_lg_do_ex4baddr153w(0) AND wire_w_lg_do_wren43w(0);
	wire_w_lg_w_lg_do_write189w190w(0) <= wire_w_lg_do_write189w(0) AND wire_w_lg_do_wren43w(0);
	wire_w_lg_w_lg_do_write53w348w(0) <= wire_w_lg_do_write53w(0) AND end_pgwr_data;
	wire_w_lg_w_lg_end_read_byte489w501w(0) <= wire_w_lg_end_read_byte489w(0) AND wire_w_lg_end_operation500w(0);
	wire_w_lg_w_lg_load_opcode160w249w(0) <= wire_w_lg_load_opcode160w(0) AND wire_w_b4addr_opcode_range248w(0);
	loop8 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode160w161w(i) <= wire_w_lg_load_opcode160w(0) AND wire_w_b4addr_opcode_range157w(i);
	END GENERATE loop8;
	wire_w_lg_w_lg_load_opcode155w247w(0) <= wire_w_lg_load_opcode155w(0) AND wire_w_exb4addr_opcode_range246w(0);
	loop9 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode155w156w(i) <= wire_w_lg_load_opcode155w(0) AND wire_w_exb4addr_opcode_range152w(i);
	END GENERATE loop9;
	wire_w_lg_w_lg_load_opcode191w263w(0) <= wire_w_lg_load_opcode191w(0) AND wire_w_write_opcode_range262w(0);
	loop10 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode191w192w(i) <= wire_w_lg_load_opcode191w(0) AND wire_w_write_opcode_range188w(i);
	END GENERATE loop10;
	wire_w_lg_w_lg_load_opcode166w167w(0) <= wire_w_lg_load_opcode166w(0) AND wire_w_lg_do_wren43w(0);
	wire_w_lg_w_lg_load_opcode171w172w(0) <= wire_w_lg_load_opcode171w(0) AND wire_w_lg_do_wren43w(0);
	wire_w_lg_w_lg_load_opcode211w271w(0) <= wire_w_lg_load_opcode211w(0) AND wire_w_fast_read_opcode_range270w(0);
	loop11 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode211w212w(i) <= wire_w_lg_load_opcode211w(0) AND wire_w_fast_read_opcode_range210w(i);
	END GENERATE loop11;
	wire_w_lg_w_lg_load_opcode214w273w(0) <= wire_w_lg_load_opcode214w(0) AND wire_w_read_opcode_range272w(0);
	loop12 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode214w215w(i) <= wire_w_lg_load_opcode214w(0) AND wire_w_read_opcode_range213w(i);
	END GENERATE loop12;
	wire_w_lg_w_lg_load_opcode194w265w(0) <= wire_w_lg_load_opcode194w(0) AND wire_w_rnvdummyclk_opcode_range264w(0);
	loop13 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode194w195w(i) <= wire_w_lg_load_opcode194w(0) AND wire_w_rnvdummyclk_opcode_range193w(i);
	END GENERATE loop13;
	wire_w_lg_w_lg_load_opcode222w277w(0) <= wire_w_lg_load_opcode222w(0) AND wire_w_rdid_opcode_range276w(0);
	loop14 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode222w223w(i) <= wire_w_lg_load_opcode222w(0) AND wire_w_rdid_opcode_range221w(i);
	END GENERATE loop14;
	wire_w_lg_w_lg_load_opcode225w279w(0) <= wire_w_lg_load_opcode225w(0) AND wire_w_rsid_opcode_range278w(0);
	loop15 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode225w226w(i) <= wire_w_lg_load_opcode225w(0) AND wire_w_rsid_opcode_range224w(i);
	END GENERATE loop15;
	wire_w_lg_w_lg_load_opcode181w186w(0) <= wire_w_lg_load_opcode181w(0) AND wire_w_lg_do_polling185w(0);
	wire_w_lg_w_lg_load_opcode181w182w(0) <= wire_w_lg_load_opcode181w(0) AND do_polling;
	wire_w_lg_w_lg_load_opcode205w206w(0) <= wire_w_lg_load_opcode205w(0) AND wire_w_lg_do_write_volatile204w(0);
	wire_w_lg_w_lg_load_opcode176w177w(0) <= wire_w_lg_load_opcode176w(0) AND wire_w_lg_do_wren43w(0);
	wire_w_lg_w_lg_load_opcode217w218w(0) <= wire_w_lg_load_opcode217w(0) AND wire_w_lg_do_wren43w(0);
	wire_w_lg_w_lg_load_opcode163w251w(0) <= wire_w_lg_load_opcode163w(0) AND wire_w_wren_opcode_range250w(0);
	loop16 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode163w164w(i) <= wire_w_lg_load_opcode163w(0) AND wire_w_wren_opcode_range162w(i);
	END GENERATE loop16;
	wire_w_lg_w_lg_load_opcode198w199w(0) <= wire_w_lg_load_opcode198w(0) AND wire_w_lg_do_read_volatile197w(0);
	wire_w_lg_w_lg_stage3_wire35w36w(0) <= wire_w_lg_stage3_wire35w(0) AND do_wait_dummyclk;
	wire_w_lg_w_lg_start_poll355w356w(0) <= wire_w_lg_start_poll355w(0) AND do_polling;
	wire_w_lg_w_lg_do_read369w370w(0) <= wire_w_lg_do_read369w(0) AND wire_w_lg_do_fast_read368w(0);
	wire_w_lg_w_lg_w_lg_w_lg_do_write62w110w111w112w(0) <= wire_w_lg_w_lg_w_lg_do_write62w110w111w(0) AND write_prot_true;
	wire_w_lg_w_lg_w_lg_do_write62w63w417w(0) <= wire_w_lg_w_lg_do_write62w63w(0) AND do_memadd;
	wire_w_lg_w_lg_do_read301w482w(0) <= wire_w_lg_do_read301w(0) AND wire_stage_cntr_w_q_range93w(0);
	wire_w_lg_w_lg_do_sec_erase44w425w(0) <= wire_w_lg_do_sec_erase44w(0) AND wire_w_lg_do_wren43w(0);
	wire_w_lg_w_lg_rden_wire421w422w(0) <= wire_w_lg_rden_wire421w(0) AND not_busy;
	wire_w_lg_addr_overdie412w(0) <= addr_overdie AND wire_w_addr_reg_overdie_range411w(0);
	loop17 : FOR i IN 0 TO 22 GENERATE 
		wire_w_lg_addr_overdie402w(i) <= addr_overdie AND wire_w_addr_reg_overdie_range401w(i);
	END GENERATE loop17;
	wire_w_lg_do_4baddr158w(0) <= do_4baddr AND wire_w_lg_do_read_stat42w(0);
	wire_w_lg_do_bulk_erase349w(0) <= do_bulk_erase AND wire_w_lg_do_read_stat42w(0);
	wire_w_lg_do_ex4baddr153w(0) <= do_ex4baddr AND wire_w_lg_do_read_stat42w(0);
	wire_w_lg_do_read_nonvolatile335w(0) <= do_read_nonvolatile AND wire_addbyte_cntr_w_q_range140w(0);
	wire_w_lg_do_write189w(0) <= do_write AND wire_w_lg_do_read_stat42w(0);
	wire_w_lg_do_write60w(0) <= do_write AND wire_w_lg_w_pagewr_buf_not_empty_range58w59w(0);
	wire_w_lg_do_write53w(0) <= do_write AND shift_pgwr_data;
	wire_w_lg_end_operation520w(0) <= end_operation AND wire_w_lg_do_read301w(0);
	wire_w_lg_end_read_byte489w(0) <= end_read_byte AND end_one_cyc_pos;
	wire_w_lg_in_operation28w(0) <= in_operation AND wire_w_lg_end_ophdly27w(0);
	wire_w_lg_load_opcode160w(0) <= load_opcode AND wire_w_lg_w_lg_do_4baddr158w159w(0);
	wire_w_lg_load_opcode155w(0) <= load_opcode AND wire_w_lg_w_lg_do_ex4baddr153w154w(0);
	wire_w_lg_load_opcode191w(0) <= load_opcode AND wire_w_lg_w_lg_do_write189w190w(0);
	wire_w_lg_load_opcode166w(0) <= load_opcode AND do_bulk_erase;
	wire_w_lg_load_opcode171w(0) <= load_opcode AND do_die_erase;
	wire_w_lg_load_opcode211w(0) <= load_opcode AND do_fast_read;
	wire_w_lg_load_opcode214w(0) <= load_opcode AND do_read;
	wire_w_lg_load_opcode194w(0) <= load_opcode AND do_read_nonvolatile;
	wire_w_lg_load_opcode222w(0) <= load_opcode AND do_read_rdid;
	wire_w_lg_load_opcode225w(0) <= load_opcode AND do_read_sid;
	wire_w_lg_load_opcode181w(0) <= load_opcode AND do_read_stat;
	wire_w_lg_load_opcode205w(0) <= load_opcode AND do_read_volatile;
	wire_w_lg_load_opcode176w(0) <= load_opcode AND do_sec_erase;
	wire_w_lg_load_opcode217w(0) <= load_opcode AND do_sec_prot;
	wire_w_lg_load_opcode163w(0) <= load_opcode AND do_wren;
	wire_w_lg_load_opcode198w(0) <= load_opcode AND do_write_volatile;
	wire_w_lg_not_busy414w(0) <= not_busy AND wire_w_addr_range413w(0);
	loop18 : FOR i IN 0 TO 22 GENERATE 
		wire_w_lg_not_busy406w(i) <= not_busy AND wire_w_addr_range405w(i);
	END GENERATE loop18;
	loop19 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_shift_opcode151w(i) <= shift_opcode AND wire_asmi_opcode_reg_w_q_range150w(i);
	END GENERATE loop19;
	wire_w_lg_stage3_wire419w(0) <= stage3_wire AND wire_w_lg_w_lg_w_lg_w_lg_do_write62w63w417w418w(0);
	wire_w_lg_stage3_wire311w(0) <= stage3_wire AND wire_w_lg_w_lg_w_lg_do_read_stat308w309w310w(0);
	wire_w_lg_stage3_wire449w(0) <= stage3_wire AND wire_w_lg_w_lg_w_lg_do_read_stat308w447w448w(0);
	wire_w_lg_stage3_wire300w(0) <= stage3_wire AND wire_w_lg_w_lg_do_read_rdid298w299w(0);
	wire_w_lg_stage3_wire45w(0) <= stage3_wire AND wire_w_lg_do_sec_erase44w(0);
	wire_w_lg_stage3_wire35w(0) <= stage3_wire AND do_fast_read;
	loop20 : FOR i IN 0 TO 22 GENERATE 
		wire_w_lg_stage3_wire404w(i) <= stage3_wire AND wire_addr_reg_w_q_range403w(i);
	END GENERATE loop20;
	wire_w_lg_stage4_wire451w(0) <= stage4_wire AND wire_w_lg_w_lg_do_read301w450w(0);
	wire_w_lg_stage4_wire302w(0) <= stage4_wire AND wire_w_lg_do_read301w(0);
	wire_w_lg_stage4_wire420w(0) <= stage4_wire AND addr_overdie;
	wire_w_lg_stage4_wire316w(0) <= stage4_wire AND do_fast_read;
	wire_w_lg_start_poll355w(0) <= start_poll AND do_read_stat;
	wire_w_lg_w_lg_do_write53w367w(0) <= NOT wire_w_lg_do_write53w(0);
	wire_w_lg_w_lg_stage4_wire316w317w(0) <= NOT wire_w_lg_stage4_wire316w(0);
	wire_w_lg_w_lg_w_lg_stage4_wire302w303w304w(0) <= NOT wire_w_lg_w_lg_stage4_wire302w303w(0);
	wire_w_lg_w_lg_w_lg_do_read_stat312w313w314w(0) <= NOT wire_w_lg_w_lg_do_read_stat312w313w(0);
	wire_w_lg_addr_overdie514w(0) <= NOT addr_overdie;
	wire_w_lg_busy_wire1w(0) <= NOT busy_wire;
	wire_w_lg_clkin_wire91w(0) <= NOT clkin_wire;
	wire_w_lg_clr_rstat_wire26w(0) <= NOT clr_rstat_wire;
	wire_w_lg_clr_sid_wire25w(0) <= NOT clr_sid_wire;
	wire_w_lg_do_fast_read368w(0) <= NOT do_fast_read;
	wire_w_lg_do_memadd434w(0) <= NOT do_memadd;
	wire_w_lg_do_polling185w(0) <= NOT do_polling;
	wire_w_lg_do_read369w(0) <= NOT do_read;
	wire_w_lg_do_read_rdid41w(0) <= NOT do_read_rdid;
	wire_w_lg_do_read_stat42w(0) <= NOT do_read_stat;
	wire_w_lg_do_read_volatile197w(0) <= NOT do_read_volatile;
	wire_w_lg_do_wren43w(0) <= NOT do_wren;
	wire_w_lg_do_write_volatile204w(0) <= NOT do_write_volatile;
	wire_w_lg_end_add_cycle73w(0) <= NOT end_add_cycle;
	wire_w_lg_end_fast_read67w(0) <= NOT end_fast_read;
	wire_w_lg_end_operation500w(0) <= NOT end_operation;
	wire_w_lg_end_ophdly27w(0) <= NOT end_ophdly;
	wire_w_lg_end_pgwr_data52w(0) <= NOT end_pgwr_data;
	wire_w_lg_end_read70w(0) <= NOT end_read;
	wire_w_lg_rden_wire516w(0) <= NOT rden_wire;
	wire_w_lg_read_rdid_wire7w(0) <= NOT read_rdid_wire;
	wire_w_lg_read_sid_wire6w(0) <= NOT read_sid_wire;
	wire_w_lg_sec_protect_wire5w(0) <= NOT sec_protect_wire;
	wire_w_lg_st_busy_wire107w(0) <= NOT st_busy_wire;
	wire_w_lg_w_pagewr_buf_not_empty_range58w59w(0) <= NOT wire_w_pagewr_buf_not_empty_range58w(0);
	wire_w_lg_w_lg_w_lg_load_opcode225w279w280w(0) <= wire_w_lg_w_lg_load_opcode225w279w(0) OR wire_w_lg_w_lg_load_opcode222w277w(0);
	loop21 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_load_opcode225w226w227w(i) <= wire_w_lg_w_lg_load_opcode225w226w(i) OR wire_w_lg_w_lg_load_opcode222w223w(i);
	END GENERATE loop21;
	wire_w_lg_w_lg_w_lg_w_lg_do_write62w63w417w418w(0) <= wire_w_lg_w_lg_w_lg_do_write62w63w417w(0) OR wire_w_lg_do_read301w(0);
	wire_w_lg_w_lg_w_lg_rden_wire421w422w423w(0) <= wire_w_lg_w_lg_rden_wire421w422w(0) OR wire_w_lg_stage4_wire420w(0);
	wire_w_lg_w_lg_not_busy414w415w(0) <= wire_w_lg_not_busy414w(0) OR wire_w_lg_addr_overdie412w(0);
	loop22 : FOR i IN 0 TO 22 GENERATE 
		wire_w_lg_w_lg_not_busy406w407w(i) <= wire_w_lg_not_busy406w(i) OR wire_w_lg_stage3_wire404w(i);
	END GENERATE loop22;
	wire_w_lg_w_lg_stage4_wire451w452w(0) <= wire_w_lg_stage4_wire451w(0) OR wire_w_lg_stage3_wire449w(0);
	wire_w_lg_w_lg_stage4_wire302w303w(0) <= wire_w_lg_stage4_wire302w(0) OR wire_w_lg_stage3_wire300w(0);
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode225w279w280w281w(0) <= wire_w_lg_w_lg_w_lg_load_opcode225w279w280w(0) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode217w218w219w275w(0);
	loop23 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_load_opcode225w226w227w228w(i) <= wire_w_lg_w_lg_w_lg_load_opcode225w226w227w(i) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode217w218w219w220w(i);
	END GENERATE loop23;
	wire_w_lg_w_lg_w_lg_w_lg_rden_wire421w422w423w424w(0) <= wire_w_lg_w_lg_w_lg_rden_wire421w422w423w(0) OR wire_w_lg_stage3_wire419w(0);
	loop24 : FOR i IN 0 TO 22 GENERATE 
		wire_w_lg_w_lg_w_lg_not_busy406w407w408w(i) <= wire_w_lg_w_lg_not_busy406w407w(i) OR wire_w_lg_addr_overdie402w(i);
	END GENERATE loop24;
	wire_w282w(0) <= wire_w_lg_w_lg_w_lg_w_lg_load_opcode225w279w280w281w(0) OR wire_w_lg_w_lg_load_opcode214w273w(0);
	loop25 : FOR i IN 0 TO 6 GENERATE 
		wire_w229w(i) <= wire_w_lg_w_lg_w_lg_w_lg_load_opcode225w226w227w228w(i) OR wire_w_lg_w_lg_load_opcode214w215w(i);
	END GENERATE loop25;
	wire_w_lg_w282w283w(0) <= wire_w282w(0) OR wire_w_lg_w_lg_load_opcode211w271w(0);
	loop26 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w229w230w(i) <= wire_w229w(i) OR wire_w_lg_w_lg_load_opcode211w212w(i);
	END GENERATE loop26;
	wire_w_lg_w_lg_w282w283w284w(0) <= wire_w_lg_w282w283w(0) OR wire_w269w(0);
	loop27 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w229w230w231w(i) <= wire_w_lg_w229w230w(i) OR wire_w209w(i);
	END GENERATE loop27;
	wire_w_lg_w_lg_w_lg_w282w283w284w285w(0) <= wire_w_lg_w_lg_w282w283w284w(0) OR wire_w267w(0);
	loop28 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w229w230w231w232w(i) <= wire_w_lg_w_lg_w229w230w231w(i) OR wire_w202w(i);
	END GENERATE loop28;
	wire_w_lg_w_lg_w_lg_w_lg_w282w283w284w285w286w(0) <= wire_w_lg_w_lg_w_lg_w282w283w284w285w(0) OR wire_w_lg_w_lg_load_opcode194w265w(0);
	loop29 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_w229w230w231w232w233w(i) <= wire_w_lg_w_lg_w_lg_w229w230w231w232w(i) OR wire_w_lg_w_lg_load_opcode194w195w(i);
	END GENERATE loop29;
	wire_w_lg_w_lg_w_lg_w_lg_w_lg_w282w283w284w285w286w287w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w282w283w284w285w286w(0) OR wire_w_lg_w_lg_load_opcode191w263w(0);
	loop30 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_w_lg_w229w230w231w232w233w234w(i) <= wire_w_lg_w_lg_w_lg_w_lg_w229w230w231w232w233w(i) OR wire_w_lg_w_lg_load_opcode191w192w(i);
	END GENERATE loop30;
	wire_w288w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w_lg_w282w283w284w285w286w287w(0) OR wire_w_lg_w_lg_w_lg_load_opcode181w186w261w(0);
	loop31 : FOR i IN 0 TO 6 GENERATE 
		wire_w235w(i) <= wire_w_lg_w_lg_w_lg_w_lg_w_lg_w229w230w231w232w233w234w(i) OR wire_w_lg_w_lg_w_lg_load_opcode181w186w187w(i);
	END GENERATE loop31;
	wire_w_lg_w288w289w(0) <= wire_w288w(0) OR wire_w_lg_w_lg_w_lg_load_opcode181w182w259w(0);
	loop32 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w235w236w(i) <= wire_w235w(i) OR wire_w_lg_w_lg_w_lg_load_opcode181w182w183w(i);
	END GENERATE loop32;
	wire_w_lg_w_lg_w288w289w290w(0) <= wire_w_lg_w288w289w(0) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode176w177w178w257w(0);
	loop33 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w235w236w237w(i) <= wire_w_lg_w235w236w(i) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode176w177w178w179w(i);
	END GENERATE loop33;
	wire_w_lg_w_lg_w_lg_w288w289w290w291w(0) <= wire_w_lg_w_lg_w288w289w290w(0) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode171w172w173w255w(0);
	loop34 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w235w236w237w238w(i) <= wire_w_lg_w_lg_w235w236w237w(i) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode171w172w173w174w(i);
	END GENERATE loop34;
	wire_w_lg_w_lg_w_lg_w_lg_w288w289w290w291w292w(0) <= wire_w_lg_w_lg_w_lg_w288w289w290w291w(0) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode166w167w168w253w(0);
	loop35 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_w235w236w237w238w239w(i) <= wire_w_lg_w_lg_w_lg_w235w236w237w238w(i) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode166w167w168w169w(i);
	END GENERATE loop35;
	wire_w_lg_w_lg_w_lg_w_lg_w_lg_w288w289w290w291w292w293w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w288w289w290w291w292w(0) OR wire_w_lg_w_lg_load_opcode163w251w(0);
	loop36 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_w_lg_w235w236w237w238w239w240w(i) <= wire_w_lg_w_lg_w_lg_w_lg_w235w236w237w238w239w(i) OR wire_w_lg_w_lg_load_opcode163w164w(i);
	END GENERATE loop36;
	wire_w294w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w_lg_w288w289w290w291w292w293w(0) OR wire_w_lg_w_lg_load_opcode160w249w(0);
	loop37 : FOR i IN 0 TO 6 GENERATE 
		wire_w241w(i) <= wire_w_lg_w_lg_w_lg_w_lg_w_lg_w235w236w237w238w239w240w(i) OR wire_w_lg_w_lg_load_opcode160w161w(i);
	END GENERATE loop37;
	wire_w_lg_w294w295w(0) <= wire_w294w(0) OR wire_w_lg_w_lg_load_opcode155w247w(0);
	loop38 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w241w242w(i) <= wire_w241w(i) OR wire_w_lg_w_lg_load_opcode155w156w(i);
	END GENERATE loop38;
	loop39 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w241w242w243w(i) <= wire_w_lg_w241w242w(i) OR wire_w_lg_shift_opcode151w(i);
	END GENERATE loop39;
	wire_w_lg_w_lg_w133w134w135w(0) <= wire_w_lg_w133w134w(0) OR do_read_nonvolatile;
	wire_w_lg_w133w134w(0) <= wire_w133w(0) OR do_fast_read;
	wire_w133w(0) <= wire_w_lg_w_lg_w_lg_w_lg_do_read_sid129w130w131w132w(0) OR do_read;
	wire_w_lg_w_lg_w_lg_w_lg_do_read301w437w438w439w(0) <= wire_w_lg_w_lg_w_lg_do_read301w437w438w(0) OR do_die_erase;
	wire_w_lg_w_lg_w_lg_w_lg_do_read_sid129w130w131w132w(0) <= wire_w_lg_w_lg_w_lg_do_read_sid129w130w131w(0) OR do_read_rdid;
	wire_w_lg_w_lg_w_lg_do_read301w437w438w(0) <= wire_w_lg_w_lg_do_read301w437w(0) OR do_sec_erase;
	wire_w_lg_w_lg_w_lg_do_read_sid129w130w131w(0) <= wire_w_lg_w_lg_do_read_sid129w130w(0) OR do_die_erase;
	wire_w_lg_w_lg_w_lg_do_read_stat308w309w310w(0) <= wire_w_lg_w_lg_do_read_stat308w309w(0) OR do_read_volatile;
	wire_w_lg_w_lg_w_lg_do_read_stat308w447w448w(0) <= wire_w_lg_w_lg_do_read_stat308w447w(0) OR do_read_nonvolatile;
	wire_w_lg_w_lg_w_lg_do_write62w110w111w(0) <= wire_w_lg_w_lg_do_write62w110w(0) OR do_die_erase;
	wire_w_lg_w_lg_do_read301w450w(0) <= wire_w_lg_do_read301w(0) OR do_read_sid;
	wire_w_lg_w_lg_do_read301w437w(0) <= wire_w_lg_do_read301w(0) OR do_write;
	wire_w_lg_w_lg_do_read_rdid298w299w(0) <= wire_w_lg_do_read_rdid298w(0) OR do_read_volatile;
	wire_w_lg_w_lg_do_read_sid129w130w(0) <= wire_w_lg_do_read_sid129w(0) OR do_sec_erase;
	wire_w_lg_w_lg_do_read_stat312w313w(0) <= wire_w_lg_do_read_stat312w(0) OR wire_w_lg_stage3_wire311w(0);
	wire_w_lg_w_lg_do_read_stat308w309w(0) <= wire_w_lg_do_read_stat308w(0) OR do_read_nonvolatile;
	wire_w_lg_w_lg_do_read_stat308w447w(0) <= wire_w_lg_do_read_stat308w(0) OR do_read_volatile;
	wire_w_lg_w_lg_do_write62w110w(0) <= wire_w_lg_do_write62w(0) OR do_bulk_erase;
	wire_w_lg_w_lg_do_write62w63w(0) <= wire_w_lg_do_write62w(0) OR do_die_erase;
	wire_w_lg_data0out_wire454w(0) <= data0out_wire OR wire_w_dataout_wire_range453w(0);
	wire_w_lg_do_4baddr351w(0) <= do_4baddr OR wire_w_lg_do_ex4baddr350w(0);
	wire_w_lg_do_ex4baddr350w(0) <= do_ex4baddr OR wire_w_lg_do_bulk_erase349w(0);
	wire_w_lg_do_read301w(0) <= do_read OR do_fast_read;
	wire_w_lg_do_read_rdid298w(0) <= do_read_rdid OR do_read_nonvolatile;
	wire_w_lg_do_read_sid129w(0) <= do_read_sid OR do_write;
	wire_w_lg_do_read_stat312w(0) <= do_read_stat OR wire_w_lg_stage4_wire302w(0);
	wire_w_lg_do_read_stat305w(0) <= do_read_stat OR wire_w_lg_w_lg_w_lg_stage4_wire302w303w304w(0);
	wire_w_lg_do_read_stat308w(0) <= do_read_stat OR do_read_rdid;
	wire_w_lg_do_sec_erase44w(0) <= do_sec_erase OR do_die_erase;
	wire_w_lg_do_wren352w(0) <= do_wren OR wire_w_lg_do_4baddr351w(0);
	wire_w_lg_do_write62w(0) <= do_write OR do_sec_erase;
	wire_w_lg_load_opcode297w(0) <= load_opcode OR shift_opcode;
	wire_w_lg_rden_wire421w(0) <= rden_wire OR wren_wire;
	add_rollover <= add_rollover_reg;
	addr_overdie <= '0';
	addr_overdie_pos <= '0';
	addr_reg_overdie <= (OTHERS => '0');
	b4addr_opcode <= (OTHERS => '0');
	berase_opcode <= (OTHERS => '0');
	busy <= busy_wire;
	busy_wire <= ((((((((((((((do_read_rdid OR do_read_sid) OR do_read) OR do_fast_read) OR do_write) OR do_sec_prot) OR do_read_stat) OR do_sec_erase) OR do_bulk_erase) OR do_die_erase) OR do_4baddr) OR do_read_volatile) OR do_fread_epcq) OR do_read_nonvolatile) OR do_ex4baddr);
	clkin_wire <= clkin;
	clr_addmsb_wire <= ((wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range93w98w429w430w(0) OR wire_w_lg_w_lg_w_lg_do_read369w370w428w(0)) OR wire_w_lg_w_lg_w_lg_w_lg_do_sec_erase44w425w426w427w(0));
	clr_endrbyte_wire <= ((((wire_w_lg_do_read301w(0) AND (NOT wire_gen_cntr_q(2))) AND wire_gen_cntr_q(1)) AND wire_gen_cntr_q(0)) OR clr_read_wire2);
	clr_read_wire <= clr_read_reg;
	clr_read_wire2 <= clr_read_reg2;
	clr_rstat_wire <= '0';
	clr_sid_wire <= '0';
	clr_write_wire2 <= '0';
	data0out_wire <= wire_sd2_data1in;
	data_valid <= data_valid_wire;
	data_valid_wire <= dvalid_reg2;
	dataoe_wire <= ( "1" & "1" & "0" & "1");
	dataout <= ( read_data_reg(7 DOWNTO 0));
	dataout_wire <= ( "0000");
	derase_opcode <= (OTHERS => '0');
	do_4baddr <= '0';
	do_bulk_erase <= '0';
	do_die_erase <= '0';
	do_ex4baddr <= '0';
	do_fast_read <= '0';
	do_fread_epcq <= '0';
	do_freadwrv_polling <= '0';
	do_memadd <= '0';
	do_polling <= ((do_write_polling OR do_sprot_polling) OR do_freadwrv_polling);
	do_read <= (((wire_w_lg_read_rdid_wire7w(0) AND wire_w_lg_read_sid_wire6w(0)) AND wire_w_lg_sec_protect_wire5w(0)) AND read_wire);
	do_read_nonvolatile <= '0';
	do_read_rdid <= '0';
	do_read_sid <= '0';
	do_read_stat <= '0';
	do_read_volatile <= '0';
	do_sec_erase <= '0';
	do_sec_prot <= '0';
	do_sprot_polling <= '0';
	do_wait_dummyclk <= '0';
	do_wren <= '0';
	do_write <= '0';
	do_write_polling <= '0';
	do_write_volatile <= '0';
	end1_cyc_gen_cntr_wire <= (wire_gen_cntr_w_lg_w_q_range103w104w(0) AND (NOT wire_gen_cntr_q(0)));
	end1_cyc_normal_in_wire <= ((((((((((wire_stage_cntr_w_lg_w_lg_w_q_range92w97w115w(0) AND (NOT wire_gen_cntr_q(2))) AND wire_gen_cntr_q(1)) AND wire_gen_cntr_q(0)) OR wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range92w97w115w116w117w(0)) OR (do_read AND end_read)) OR (do_fast_read AND end_fast_read)) OR wire_w_lg_w_lg_w_lg_w_lg_do_write62w110w111w112w(0)) OR wire_w_lg_do_write60w(0)) OR ((do_read_stat AND start_poll) AND wire_w_lg_st_busy_wire107w(0))) OR (do_read_rdid AND end_op_wire));
	end1_cyc_reg_in_wire <= end1_cyc_normal_in_wire;
	end_add_cycle <= wire_mux211_dataout;
	end_add_cycle_mux_datab_wire <= (wire_addbyte_cntr_q(2) AND wire_addbyte_cntr_q(1));
	end_fast_read <= end_read_reg;
	end_one_cyc_pos <= end1_cyc_reg2;
	end_one_cycle <= end1_cyc_reg;
	end_op_wire <= (((((((((((wire_stage_cntr_w_lg_w_q_range93w98w(0) AND ((wire_w_lg_w_lg_w_lg_w_lg_do_read369w370w371w372w(0) OR (do_read AND end_read)) OR (do_fast_read AND end_fast_read))) OR (wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range93w96w364w365w(0) AND wire_w_lg_do_polling185w(0))) OR ((((((do_read_rdid AND end_one_cyc_pos) AND wire_stage_cntr_q(1)) AND wire_stage_cntr_q(0)) AND wire_addbyte_cntr_q(2)) AND wire_addbyte_cntr_q(1)) AND wire_addbyte_cntr_w_lg_w_q_range143w144w(0))) OR (wire_w_lg_w_lg_start_poll355w356w(0) AND wire_w_lg_st_busy_wire107w(0))) OR wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range93w94w95w353w354w(0)) OR wire_w_lg_w_lg_w_lg_w_lg_do_write62w110w111w112w(0)) OR wire_w_lg_w_lg_do_write53w348w(0)) OR wire_w_lg_do_write60w(0)) OR wire_stage_cntr_w347w(0)) OR wire_stage_cntr_w_lg_w342w343w(0)) OR (wire_stage_cntr_w_lg_w_lg_w_q_range93w96w337w(0) AND ((do_write_volatile OR do_read_volatile) OR wire_w_lg_do_read_nonvolatile335w(0))));
	end_operation <= end_op_reg;
	end_ophdly <= end_op_hdlyreg;
	end_pgwr_data <= '0';
	end_read <= end_read_reg;
	end_read_byte <= (end_rbyte_reg AND wire_w_lg_addr_overdie514w(0));
	exb4addr_opcode <= (OTHERS => '0');
	fast_read_opcode <= (OTHERS => '0');
	freadwrv_sdoin <= '0';
	in_operation <= busy_wire;
	load_opcode <= ((((wire_stage_cntr_w_lg_w_q_range93w94w(0) AND wire_stage_cntr_w_lg_w_q_range92w97w(0)) AND (NOT wire_gen_cntr_q(2))) AND wire_gen_cntr_w_lg_w_q_range101w102w(0)) AND wire_gen_cntr_q(0));
	memadd_sdoin <= add_msb_reg;
	ncs_reg_ena_wire <= (((wire_stage_cntr_w_lg_w_lg_w_q_range93w94w95w(0) AND end_one_cyc_pos) OR addr_overdie_pos) OR end_operation);
	not_busy <= busy_det_reg;
	oe_wire <= '0';
	pagewr_buf_not_empty <= ( "1");
	rden_wire <= rden;
	rdid_opcode <= (OTHERS => '0');
	rdummyclk_opcode <= (OTHERS => '0');
	read_address <= ( read_add_reg(23 DOWNTO 0));
	read_data_reg_in_wire <= ( read_dout_reg(7 DOWNTO 0));
	read_opcode <= "00000011";
	read_rdid_wire <= '0';
	read_sid_wire <= '0';
	read_wire <= read_reg;
	rflagstat_opcode <= (OTHERS => '0');
	rnvdummyclk_opcode <= (OTHERS => '0');
	rsid_opcode <= (OTHERS => '0');
	rsid_sdoin <= '0';
	rstat_opcode <= (OTHERS => '0');
	scein_wire <= wire_ncs_reg_w_lg_q390w(0);
	sdoin_wire <= to_sdoin_wire;
	sec_protect_wire <= '0';
	secprot_opcode <= (OTHERS => '0');
	secprot_sdoin <= '0';
	serase_opcode <= (OTHERS => '0');
	shift_opcode <= shift_op_reg;
	shift_opdata <= stage2_wire;
	shift_pgwr_data <= '0';
	st_busy_wire <= '0';
	stage2_wire <= stage2_reg;
	stage3_wire <= stage3_reg;
	stage4_wire <= stage4_reg;
	start_frpoll <= '0';
	start_poll <= ((start_wrpoll OR start_sppoll) OR start_frpoll);
	start_sppoll <= '0';
	start_wrpoll <= '0';
	to_sdoin_wire <= ((((((shift_opdata AND asmi_opcode_reg(7)) OR rsid_sdoin) OR memadd_sdoin) OR write_sdoin) OR secprot_sdoin) OR freadwrv_sdoin);
	wren_opcode <= (OTHERS => '0');
	wren_wire <= '1';
	write_opcode <= (OTHERS => '0');
	write_prot_true <= '0';
	write_sdoin <= '0';
	wrvolatile_opcode <= (OTHERS => '0');
	wire_w_addr_range413w(0) <= addr(0);
	wire_w_addr_range405w <= addr(23 DOWNTO 1);
	wire_w_addr_reg_overdie_range411w(0) <= addr_reg_overdie(0);
	wire_w_addr_reg_overdie_range401w <= addr_reg_overdie(23 DOWNTO 1);
	wire_w_b4addr_opcode_range248w(0) <= b4addr_opcode(0);
	wire_w_b4addr_opcode_range157w <= b4addr_opcode(7 DOWNTO 1);
	wire_w_berase_opcode_range252w(0) <= berase_opcode(0);
	wire_w_berase_opcode_range165w <= berase_opcode(7 DOWNTO 1);
	wire_w_dataout_wire_range453w(0) <= dataout_wire(1);
	wire_w_derase_opcode_range254w(0) <= derase_opcode(0);
	wire_w_derase_opcode_range170w <= derase_opcode(7 DOWNTO 1);
	wire_w_exb4addr_opcode_range246w(0) <= exb4addr_opcode(0);
	wire_w_exb4addr_opcode_range152w <= exb4addr_opcode(7 DOWNTO 1);
	wire_w_fast_read_opcode_range270w(0) <= fast_read_opcode(0);
	wire_w_fast_read_opcode_range210w <= fast_read_opcode(7 DOWNTO 1);
	wire_w_pagewr_buf_not_empty_range58w(0) <= pagewr_buf_not_empty(0);
	wire_w_rdid_opcode_range276w(0) <= rdid_opcode(0);
	wire_w_rdid_opcode_range221w <= rdid_opcode(7 DOWNTO 1);
	wire_w_rdummyclk_opcode_range268w(0) <= rdummyclk_opcode(0);
	wire_w_rdummyclk_opcode_range203w <= rdummyclk_opcode(7 DOWNTO 1);
	wire_w_read_opcode_range272w(0) <= read_opcode(0);
	wire_w_read_opcode_range213w <= read_opcode(7 DOWNTO 1);
	wire_w_rflagstat_opcode_range258w(0) <= rflagstat_opcode(0);
	wire_w_rflagstat_opcode_range180w <= rflagstat_opcode(7 DOWNTO 1);
	wire_w_rnvdummyclk_opcode_range264w(0) <= rnvdummyclk_opcode(0);
	wire_w_rnvdummyclk_opcode_range193w <= rnvdummyclk_opcode(7 DOWNTO 1);
	wire_w_rsid_opcode_range278w(0) <= rsid_opcode(0);
	wire_w_rsid_opcode_range224w <= rsid_opcode(7 DOWNTO 1);
	wire_w_rstat_opcode_range260w(0) <= rstat_opcode(0);
	wire_w_rstat_opcode_range184w <= rstat_opcode(7 DOWNTO 1);
	wire_w_secprot_opcode_range274w(0) <= secprot_opcode(0);
	wire_w_secprot_opcode_range216w <= secprot_opcode(7 DOWNTO 1);
	wire_w_serase_opcode_range256w(0) <= serase_opcode(0);
	wire_w_serase_opcode_range175w <= serase_opcode(7 DOWNTO 1);
	wire_w_wren_opcode_range250w(0) <= wren_opcode(0);
	wire_w_wren_opcode_range162w <= wren_opcode(7 DOWNTO 1);
	wire_w_write_opcode_range262w(0) <= write_opcode(0);
	wire_w_write_opcode_range188w <= write_opcode(7 DOWNTO 1);
	wire_w_wrvolatile_opcode_range266w(0) <= wrvolatile_opcode(0);
	wire_w_wrvolatile_opcode_range196w <= wrvolatile_opcode(7 DOWNTO 1);
	wire_addbyte_cntr_w_lg_w_q_range140w145w(0) <= wire_addbyte_cntr_w_q_range140w(0) AND wire_addbyte_cntr_w_lg_w_q_range143w144w(0);
	wire_addbyte_cntr_w_lg_w_q_range143w144w(0) <= NOT wire_addbyte_cntr_w_q_range143w(0);
	wire_addbyte_cntr_clk_en <= wire_stage_cntr_w139w(0);
	wire_stage_cntr_w139w(0) <= ((wire_stage_cntr_w_lg_w_lg_w_q_range93w96w136w(0) AND wire_w_lg_w_lg_w133w134w135w(0)) OR addr_overdie) OR end_operation;
	wire_addbyte_cntr_clock <= wire_w_lg_clkin_wire91w(0);
	wire_addbyte_cntr_sclr <= wire_w_lg_end_operation90w(0);
	wire_w_lg_end_operation90w(0) <= end_operation OR addr_overdie;
	wire_addbyte_cntr_w_q_range143w(0) <= wire_addbyte_cntr_q(0);
	wire_addbyte_cntr_w_q_range140w(0) <= wire_addbyte_cntr_q(1);
	addbyte_cntr :  a_graycounter
	  GENERIC MAP (
		WIDTH => 3
	  )
	  PORT MAP ( 
		aclr => reset,
		clk_en => wire_addbyte_cntr_clk_en,
		clock => wire_addbyte_cntr_clock,
		q => wire_addbyte_cntr_q,
		sclr => wire_addbyte_cntr_sclr
	  );
	wire_gen_cntr_w_lg_w_q_range103w104w(0) <= wire_gen_cntr_w_q_range103w(0) AND wire_gen_cntr_w_lg_w_q_range101w102w(0);
	wire_gen_cntr_w_lg_w_q_range101w102w(0) <= NOT wire_gen_cntr_w_q_range101w(0);
	wire_gen_cntr_clk_en <= wire_w32w(0);
	wire_w32w(0) <= (((wire_w_lg_in_operation28w(0) AND wire_w_lg_clr_rstat_wire26w(0)) AND wire_w_lg_clr_sid_wire25w(0)) OR do_wait_dummyclk) OR addr_overdie;
	wire_gen_cntr_sclr <= wire_w_lg_w_lg_end1_cyc_reg_in_wire33w34w(0);
	wire_w_lg_w_lg_end1_cyc_reg_in_wire33w34w(0) <= (end1_cyc_reg_in_wire OR addr_overdie) OR do_wait_dummyclk;
	wire_gen_cntr_w_q_range101w(0) <= wire_gen_cntr_q(1);
	wire_gen_cntr_w_q_range103w(0) <= wire_gen_cntr_q(2);
	gen_cntr :  a_graycounter
	  GENERIC MAP (
		WIDTH => 3
	  )
	  PORT MAP ( 
		aclr => reset,
		clk_en => wire_gen_cntr_clk_en,
		clock => clkin_wire,
		q => wire_gen_cntr_q,
		sclr => wire_gen_cntr_sclr
	  );
	wire_stage_cntr_w_lg_w342w343w(0) <= wire_stage_cntr_w342w(0) AND end_one_cycle;
	wire_stage_cntr_w342w(0) <= wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range93w96w339w340w341w(0) AND end_add_cycle;
	wire_stage_cntr_w347w(0) <= wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range93w96w344w345w346w(0) AND end_one_cycle;
	wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range93w96w339w340w341w(0) <= wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range93w96w339w340w(0) AND wire_w_lg_do_read_stat42w(0);
	wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range93w96w344w345w346w(0) <= wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range93w96w344w345w(0) AND wire_w_lg_do_read_stat42w(0);
	wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range93w94w95w353w354w(0) <= wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range93w94w95w353w(0) AND end_one_cycle;
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range93w98w429w430w(0) <= wire_stage_cntr_w_lg_w_lg_w_q_range93w98w429w(0) AND end_one_cyc_pos;
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range93w96w339w340w(0) <= wire_stage_cntr_w_lg_w_lg_w_q_range93w96w339w(0) AND wire_w_lg_do_wren43w(0);
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range93w96w364w365w(0) <= wire_stage_cntr_w_lg_w_lg_w_q_range93w96w364w(0) AND end_one_cycle;
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range93w96w344w345w(0) <= wire_stage_cntr_w_lg_w_lg_w_q_range93w96w344w(0) AND wire_w_lg_do_wren43w(0);
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range93w94w95w353w(0) <= wire_stage_cntr_w_lg_w_lg_w_q_range93w94w95w(0) AND wire_w_lg_do_wren352w(0);
	wire_stage_cntr_w_lg_w_lg_w_q_range93w98w429w(0) <= wire_stage_cntr_w_lg_w_q_range93w98w(0) AND end_add_cycle;
	wire_stage_cntr_w_lg_w_lg_w_q_range93w96w339w(0) <= wire_stage_cntr_w_lg_w_q_range93w96w(0) AND wire_w_lg_do_sec_erase44w(0);
	wire_stage_cntr_w_lg_w_lg_w_q_range93w96w364w(0) <= wire_stage_cntr_w_lg_w_q_range93w96w(0) AND do_read_stat;
	wire_stage_cntr_w_lg_w_lg_w_q_range93w96w344w(0) <= wire_stage_cntr_w_lg_w_q_range93w96w(0) AND do_sec_prot;
	wire_stage_cntr_w_lg_w_lg_w_q_range93w96w136w(0) <= wire_stage_cntr_w_lg_w_q_range93w96w(0) AND end_one_cyc_pos;
	wire_stage_cntr_w_lg_w_lg_w_q_range93w96w337w(0) <= wire_stage_cntr_w_lg_w_q_range93w96w(0) AND end_one_cycle;
	wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range92w97w115w116w117w(0) <= wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range92w97w115w116w(0) AND end1_cyc_gen_cntr_wire;
	wire_stage_cntr_w_lg_w_lg_w_q_range92w97w115w(0) <= wire_stage_cntr_w_lg_w_q_range92w97w(0) AND wire_stage_cntr_w_lg_w_q_range93w94w(0);
	wire_stage_cntr_w_lg_w_lg_w_q_range93w94w95w(0) <= wire_stage_cntr_w_lg_w_q_range93w94w(0) AND wire_stage_cntr_w_q_range92w(0);
	wire_stage_cntr_w_lg_w_q_range93w98w(0) <= wire_stage_cntr_w_q_range93w(0) AND wire_stage_cntr_w_lg_w_q_range92w97w(0);
	wire_stage_cntr_w_lg_w_q_range93w96w(0) <= wire_stage_cntr_w_q_range93w(0) AND wire_stage_cntr_w_q_range92w(0);
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range92w97w115w116w(0) <= NOT wire_stage_cntr_w_lg_w_lg_w_q_range92w97w115w(0);
	wire_stage_cntr_w_lg_w_q_range92w97w(0) <= NOT wire_stage_cntr_w_q_range92w(0);
	wire_stage_cntr_w_lg_w_q_range93w94w(0) <= NOT wire_stage_cntr_w_q_range93w(0);
	wire_stage_cntr_clk_en <= wire_w_lg_w_lg_w_lg_w86w87w88w89w(0);
	wire_w_lg_w_lg_w_lg_w86w87w88w89w(0) <= (((((((((((((in_operation AND end_one_cycle) AND (NOT (stage3_wire AND wire_w_lg_end_add_cycle73w(0)))) AND (NOT (stage4_wire AND wire_w_lg_end_read70w(0)))) AND (NOT (stage4_wire AND wire_w_lg_end_fast_read67w(0)))) AND (NOT ((wire_w_lg_w_lg_do_write62w63w(0) OR do_bulk_erase) AND write_prot_true))) AND (NOT wire_w_lg_do_write60w(0))) AND (NOT (stage3_wire AND st_busy_wire))) AND (NOT (wire_w_lg_do_write53w(0) AND wire_w_lg_end_pgwr_data52w(0)))) AND (NOT (stage2_wire AND do_wren))) AND (NOT (((wire_w_lg_stage3_wire45w(0) AND wire_w_lg_do_wren43w(0)) AND wire_w_lg_do_read_stat42w(0)) AND wire_w_lg_do_read_rdid41w(0)))) AND (NOT (stage3_wire AND ((do_write_volatile OR do_read_volatile) OR do_read_nonvolatile)))) OR wire_w_lg_w_lg_stage3_wire35w36w(0)) OR addr_overdie) OR end_ophdly;
	wire_stage_cntr_sclr <= wire_w_lg_end_operation90w(0);
	wire_stage_cntr_w_q_range92w(0) <= wire_stage_cntr_q(0);
	wire_stage_cntr_w_q_range93w(0) <= wire_stage_cntr_q(1);
	stage_cntr :  a_graycounter
	  GENERIC MAP (
		WIDTH => 2
	  )
	  PORT MAP ( 
		aclr => reset,
		clk_en => wire_stage_cntr_clk_en,
		clock => clkin_wire,
		q => wire_stage_cntr_q,
		sclr => wire_stage_cntr_sclr
	  );
	sd2 :  cyclonev_asmiblock
	  GENERIC MAP (
		enable_sim => "false"
	  )
	  PORT MAP ( 
		data0oe => dataoe_wire(0),
		data0out => sdoin_wire,
		data1in => wire_sd2_data1in,
		data1oe => dataoe_wire(1),
		data2oe => dataoe_wire(2),
		data2out => wire_vcc,
		data3oe => dataoe_wire(3),
		data3out => wire_vcc,
		dclk => clkin_wire,
		oe => oe_wire,
		sce => scein_wire
	  );
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN add_msb_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_add_msb_reg_ena = '1') THEN 
				IF (clr_addmsb_wire = '1') THEN add_msb_reg <= '0';
				ELSE add_msb_reg <= addr_reg(23);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_add_msb_reg_ena <= ((((wire_w_lg_w_lg_w_lg_w_lg_do_read301w437w438w439w(0) AND (NOT (wire_w_lg_w_lg_do_write62w63w(0) AND wire_w_lg_do_memadd434w(0)))) AND wire_stage_cntr_q(1)) AND wire_stage_cntr_q(0)) OR clr_addmsb_wire);
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN add_rollover_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN add_rollover_reg <= (wire_read_add_cntr_q(23) OR clr_read_wire2);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(0) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(0) = '1') THEN addr_reg(0) <= wire_addr_reg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(1) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(1) = '1') THEN addr_reg(1) <= wire_addr_reg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(2) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(2) = '1') THEN addr_reg(2) <= wire_addr_reg_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(3) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(3) = '1') THEN addr_reg(3) <= wire_addr_reg_d(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(4) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(4) = '1') THEN addr_reg(4) <= wire_addr_reg_d(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(5) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(5) = '1') THEN addr_reg(5) <= wire_addr_reg_d(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(6) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(6) = '1') THEN addr_reg(6) <= wire_addr_reg_d(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(7) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(7) = '1') THEN addr_reg(7) <= wire_addr_reg_d(7);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(8) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(8) = '1') THEN addr_reg(8) <= wire_addr_reg_d(8);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(9) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(9) = '1') THEN addr_reg(9) <= wire_addr_reg_d(9);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(10) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(10) = '1') THEN addr_reg(10) <= wire_addr_reg_d(10);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(11) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(11) = '1') THEN addr_reg(11) <= wire_addr_reg_d(11);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(12) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(12) = '1') THEN addr_reg(12) <= wire_addr_reg_d(12);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(13) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(13) = '1') THEN addr_reg(13) <= wire_addr_reg_d(13);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(14) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(14) = '1') THEN addr_reg(14) <= wire_addr_reg_d(14);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(15) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(15) = '1') THEN addr_reg(15) <= wire_addr_reg_d(15);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(16) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(16) = '1') THEN addr_reg(16) <= wire_addr_reg_d(16);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(17) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(17) = '1') THEN addr_reg(17) <= wire_addr_reg_d(17);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(18) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(18) = '1') THEN addr_reg(18) <= wire_addr_reg_d(18);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(19) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(19) = '1') THEN addr_reg(19) <= wire_addr_reg_d(19);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(20) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(20) = '1') THEN addr_reg(20) <= wire_addr_reg_d(20);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(21) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(21) = '1') THEN addr_reg(21) <= wire_addr_reg_d(21);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(22) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(22) = '1') THEN addr_reg(22) <= wire_addr_reg_d(22);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(23) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(23) = '1') THEN addr_reg(23) <= wire_addr_reg_d(23);
			END IF;
		END IF;
	END PROCESS;
	wire_addr_reg_d <= ( wire_w_lg_w_lg_w_lg_not_busy406w407w408w & wire_w_lg_w_lg_not_busy414w415w);
	loop40 : FOR i IN 0 TO 23 GENERATE
		wire_addr_reg_ena(i) <= wire_w_lg_w_lg_w_lg_w_lg_rden_wire421w422w423w424w(0);
	END GENERATE loop40;
	wire_addr_reg_w_q_range403w <= addr_reg(22 DOWNTO 0);
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN asmi_opcode_reg(0) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(0) = '1') THEN asmi_opcode_reg(0) <= wire_asmi_opcode_reg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN asmi_opcode_reg(1) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(1) = '1') THEN asmi_opcode_reg(1) <= wire_asmi_opcode_reg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN asmi_opcode_reg(2) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(2) = '1') THEN asmi_opcode_reg(2) <= wire_asmi_opcode_reg_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN asmi_opcode_reg(3) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(3) = '1') THEN asmi_opcode_reg(3) <= wire_asmi_opcode_reg_d(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN asmi_opcode_reg(4) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(4) = '1') THEN asmi_opcode_reg(4) <= wire_asmi_opcode_reg_d(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN asmi_opcode_reg(5) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(5) = '1') THEN asmi_opcode_reg(5) <= wire_asmi_opcode_reg_d(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN asmi_opcode_reg(6) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(6) = '1') THEN asmi_opcode_reg(6) <= wire_asmi_opcode_reg_d(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN asmi_opcode_reg(7) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(7) = '1') THEN asmi_opcode_reg(7) <= wire_asmi_opcode_reg_d(7);
			END IF;
		END IF;
	END PROCESS;
	wire_asmi_opcode_reg_d <= ( wire_w_lg_w_lg_w241w242w243w & wire_w_lg_w294w295w);
	loop41 : FOR i IN 0 TO 7 GENERATE
		wire_asmi_opcode_reg_ena(i) <= wire_w_lg_load_opcode297w(0);
	END GENERATE loop41;
	wire_asmi_opcode_reg_w_q_range150w <= asmi_opcode_reg(6 DOWNTO 0);
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN busy_det_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN busy_det_reg <= wire_w_lg_busy_wire1w(0);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN clr_read_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN clr_read_reg <= ((do_read_sid OR do_sec_prot) OR wire_w_lg_end_operation520w(0));
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN clr_read_reg2 <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN clr_read_reg2 <= clr_read_reg;
		END IF;
	END PROCESS;
	dffe3 <= '0';
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN dvalid_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_dvalid_reg_ena = '1') THEN 
				IF (wire_dvalid_reg_sclr = '1') THEN dvalid_reg <= '0';
				ELSE dvalid_reg <= wire_w_lg_end_read_byte489w(0);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_dvalid_reg_ena <= wire_w_lg_do_read301w(0);
	wire_dvalid_reg_sclr <= (end_op_wire OR end_operation);
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN dvalid_reg2 <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN dvalid_reg2 <= dvalid_reg;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN end1_cyc_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN end1_cyc_reg <= end1_cyc_reg_in_wire;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN end1_cyc_reg2 <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN end1_cyc_reg2 <= end_one_cycle;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN end_op_hdlyreg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN end_op_hdlyreg <= end_operation;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN end_op_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN end_op_reg <= end_op_wire;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN end_rbyte_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_end_rbyte_reg_ena = '1') THEN 
				IF (wire_end_rbyte_reg_sclr = '1') THEN end_rbyte_reg <= '0';
				ELSE end_rbyte_reg <= wire_w_lg_w_lg_w_lg_do_read301w482w483w(0);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_end_rbyte_reg_ena <= ((wire_gen_cntr_w_lg_w_q_range103w104w(0) AND wire_gen_cntr_q(0)) OR clr_endrbyte_wire);
	wire_end_rbyte_reg_sclr <= (clr_endrbyte_wire OR addr_overdie);
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN end_read_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN end_read_reg <= (((wire_w_lg_rden_wire516w(0) AND wire_w_lg_do_read301w(0)) AND data_valid_wire) AND end_read_byte);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN ncs_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (ncs_reg_ena_wire = '1') THEN 
				IF (wire_ncs_reg_sclr = '1') THEN ncs_reg <= '0';
				ELSE ncs_reg <= '1';
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_ncs_reg_sclr <= (end_operation OR addr_overdie_pos);
	wire_ncs_reg_w_lg_q390w(0) <= NOT ncs_reg;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(0) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(0) = '1') THEN read_add_reg(0) <= wire_read_add_reg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(1) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(1) = '1') THEN read_add_reg(1) <= wire_read_add_reg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(2) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(2) = '1') THEN read_add_reg(2) <= wire_read_add_reg_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(3) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(3) = '1') THEN read_add_reg(3) <= wire_read_add_reg_d(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(4) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(4) = '1') THEN read_add_reg(4) <= wire_read_add_reg_d(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(5) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(5) = '1') THEN read_add_reg(5) <= wire_read_add_reg_d(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(6) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(6) = '1') THEN read_add_reg(6) <= wire_read_add_reg_d(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(7) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(7) = '1') THEN read_add_reg(7) <= wire_read_add_reg_d(7);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(8) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(8) = '1') THEN read_add_reg(8) <= wire_read_add_reg_d(8);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(9) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(9) = '1') THEN read_add_reg(9) <= wire_read_add_reg_d(9);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(10) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(10) = '1') THEN read_add_reg(10) <= wire_read_add_reg_d(10);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(11) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(11) = '1') THEN read_add_reg(11) <= wire_read_add_reg_d(11);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(12) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(12) = '1') THEN read_add_reg(12) <= wire_read_add_reg_d(12);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(13) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(13) = '1') THEN read_add_reg(13) <= wire_read_add_reg_d(13);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(14) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(14) = '1') THEN read_add_reg(14) <= wire_read_add_reg_d(14);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(15) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(15) = '1') THEN read_add_reg(15) <= wire_read_add_reg_d(15);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(16) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(16) = '1') THEN read_add_reg(16) <= wire_read_add_reg_d(16);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(17) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(17) = '1') THEN read_add_reg(17) <= wire_read_add_reg_d(17);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(18) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(18) = '1') THEN read_add_reg(18) <= wire_read_add_reg_d(18);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(19) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(19) = '1') THEN read_add_reg(19) <= wire_read_add_reg_d(19);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(20) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(20) = '1') THEN read_add_reg(20) <= wire_read_add_reg_d(20);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(21) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(21) = '1') THEN read_add_reg(21) <= wire_read_add_reg_d(21);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(22) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(22) = '1') THEN read_add_reg(22) <= wire_read_add_reg_d(22);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(23) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(23) = '1') THEN read_add_reg(23) <= wire_read_add_reg_d(23);
			END IF;
		END IF;
	END PROCESS;
	wire_read_add_reg_d <= ( wire_read_add_cntr_q(23 DOWNTO 0));
	loop42 : FOR i IN 0 TO 23 GENERATE
		wire_read_add_reg_ena(i) <= wire_w_lg_w_lg_end_read_byte489w501w(0);
	END GENERATE loop42;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_data_reg(0) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(0) = '1') THEN read_data_reg(0) <= wire_read_data_reg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_data_reg(1) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(1) = '1') THEN read_data_reg(1) <= wire_read_data_reg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_data_reg(2) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(2) = '1') THEN read_data_reg(2) <= wire_read_data_reg_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_data_reg(3) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(3) = '1') THEN read_data_reg(3) <= wire_read_data_reg_d(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_data_reg(4) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(4) = '1') THEN read_data_reg(4) <= wire_read_data_reg_d(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_data_reg(5) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(5) = '1') THEN read_data_reg(5) <= wire_read_data_reg_d(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_data_reg(6) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(6) = '1') THEN read_data_reg(6) <= wire_read_data_reg_d(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_data_reg(7) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(7) = '1') THEN read_data_reg(7) <= wire_read_data_reg_d(7);
			END IF;
		END IF;
	END PROCESS;
	wire_read_data_reg_d <= ( read_data_reg_in_wire(7 DOWNTO 0));
	loop43 : FOR i IN 0 TO 7 GENERATE
		wire_read_data_reg_ena(i) <= wire_w485w(0);
	END GENERATE loop43;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_dout_reg(0) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(0) = '1') THEN read_dout_reg(0) <= wire_read_dout_reg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_dout_reg(1) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(1) = '1') THEN read_dout_reg(1) <= wire_read_dout_reg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_dout_reg(2) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(2) = '1') THEN read_dout_reg(2) <= wire_read_dout_reg_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_dout_reg(3) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(3) = '1') THEN read_dout_reg(3) <= wire_read_dout_reg_d(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_dout_reg(4) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(4) = '1') THEN read_dout_reg(4) <= wire_read_dout_reg_d(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_dout_reg(5) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(5) = '1') THEN read_dout_reg(5) <= wire_read_dout_reg_d(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_dout_reg(6) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(6) = '1') THEN read_dout_reg(6) <= wire_read_dout_reg_d(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_dout_reg(7) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(7) = '1') THEN read_dout_reg(7) <= wire_read_dout_reg_d(7);
			END IF;
		END IF;
	END PROCESS;
	wire_read_dout_reg_d <= ( read_dout_reg(6 DOWNTO 0) & wire_w_lg_data0out_wire454w);
	loop44 : FOR i IN 0 TO 7 GENERATE
		wire_read_dout_reg_ena(i) <= wire_w_lg_w_lg_stage4_wire451w452w(0);
	END GENERATE loop44;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_reg_ena = '1') THEN 
				IF (clr_read_wire = '1') THEN read_reg <= '0';
				ELSE read_reg <= read;
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_read_reg_ena <= ((wire_w_lg_busy_wire1w(0) AND rden_wire) OR clr_read_wire);
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN shift_op_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN shift_op_reg <= wire_stage_cntr_w_lg_w_lg_w_q_range93w94w95w(0);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN stage2_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN stage2_reg <= wire_stage_cntr_w_lg_w_lg_w_q_range93w94w95w(0);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN stage3_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN stage3_reg <= wire_stage_cntr_w_lg_w_q_range93w96w(0);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN stage4_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN stage4_reg <= wire_stage_cntr_w_lg_w_q_range93w98w(0);
		END IF;
	END PROCESS;
	wire_read_add_cntr_clk_en <= wire_w_lg_w_lg_w_lg_rden_wire491w492w493w(0);
	wire_w_lg_w_lg_w_lg_rden_wire491w492w493w(0) <= ((rden_wire AND not_busy) OR data_valid_wire) OR add_rollover;
	wire_read_add_cntr_data <= ( "0" & addr(23 DOWNTO 0));
	wire_read_add_cntr_sload <= wire_w_lg_rden_wire491w(0);
	wire_w_lg_rden_wire491w(0) <= rden_wire AND not_busy;
	read_add_cntr :  lpm_counter
	  GENERIC MAP (
		lpm_direction => "UP",
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 25
	  )
	  PORT MAP ( 
		aclr => reset,
		clk_en => wire_read_add_cntr_clk_en,
		clock => clkin_wire,
		data => wire_read_add_cntr_data,
		q => wire_read_add_cntr_q,
		sclr => add_rollover,
		sload => wire_read_add_cntr_sload
	  );
	wire_mux211_dataout <= end_add_cycle_mux_datab_wire WHEN do_fast_read = '1'  ELSE wire_addbyte_cntr_w_lg_w_q_range140w145w(0);

 END RTL; --asmicont_altasmi_parallel_ehl2
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY asmicont IS
	PORT
	(
		addr		: IN STD_LOGIC_VECTOR (23 DOWNTO 0);
		clkin		: IN STD_LOGIC ;
		rden		: IN STD_LOGIC ;
		read		: IN STD_LOGIC ;
		reset		: IN STD_LOGIC ;
		busy		: OUT STD_LOGIC ;
		data_valid		: OUT STD_LOGIC ;
		dataout		: OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
		read_address		: OUT STD_LOGIC_VECTOR (23 DOWNTO 0)
	);
END asmicont;


ARCHITECTURE RTL OF asmicont IS

	ATTRIBUTE synthesis_clearbox: natural;
	ATTRIBUTE synthesis_clearbox OF RTL: ARCHITECTURE IS 2;
	ATTRIBUTE clearbox_macroname: string;
	ATTRIBUTE clearbox_macroname OF RTL: ARCHITECTURE IS "ALTASMI_PARALLEL";
	ATTRIBUTE clearbox_defparam: string;
	ATTRIBUTE clearbox_defparam OF RTL: ARCHITECTURE IS "data_width=STANDARD;enable_sim=FALSE;epcs_type=EPCS64;flash_rstpin=FALSE;intended_device_family=Cyclone V;lpm_hint=UNUSED;lpm_type=altasmi_parallel;page_size=1;port_bulk_erase=PORT_UNUSED;port_die_erase=PORT_UNUSED;port_en4b_addr=PORT_UNUSED;port_ex4b_addr=PORT_UNUSED;port_fast_read=PORT_UNUSED;port_illegal_erase=PORT_UNUSED;port_illegal_write=PORT_UNUSED;port_rdid_out=PORT_UNUSED;port_read_address=PORT_USED;port_read_dummyclk=PORT_UNUSED;port_read_rdid=PORT_UNUSED;port_read_sid=PORT_UNUSED;port_read_status=PORT_UNUSED;port_sector_erase=PORT_UNUSED;port_sector_protect=PORT_UNUSED;port_shift_bytes=PORT_UNUSED;port_wren=PORT_UNUSED;port_write=PORT_UNUSED;use_asmiblock=ON;use_eab=ON;write_dummy_clk=0;";
	SIGNAL sub_wire0	: STD_LOGIC ;
	SIGNAL sub_wire1	: STD_LOGIC ;
	SIGNAL sub_wire2	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire3	: STD_LOGIC_VECTOR (23 DOWNTO 0);



	COMPONENT asmicont_altasmi_parallel_ehl2
	PORT (
			addr	: IN STD_LOGIC_VECTOR (23 DOWNTO 0);
			clkin	: IN STD_LOGIC ;
			rden	: IN STD_LOGIC ;
			read	: IN STD_LOGIC ;
			reset	: IN STD_LOGIC ;
			busy	: OUT STD_LOGIC ;
			data_valid	: OUT STD_LOGIC ;
			dataout	: OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
			read_address	: OUT STD_LOGIC_VECTOR (23 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	busy    <= sub_wire0;
	data_valid    <= sub_wire1;
	dataout    <= sub_wire2(7 DOWNTO 0);
	read_address    <= sub_wire3(23 DOWNTO 0);

	asmicont_altasmi_parallel_ehl2_component : asmicont_altasmi_parallel_ehl2
	PORT MAP (
		addr => addr,
		clkin => clkin,
		rden => rden,
		read => read,
		reset => reset,
		busy => sub_wire0,
		data_valid => sub_wire1,
		dataout => sub_wire2,
		read_address => sub_wire3
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
-- Retrieval info: CONSTANT: DATA_WIDTH STRING "STANDARD"
-- Retrieval info: CONSTANT: ENABLE_SIM STRING "FALSE"
-- Retrieval info: CONSTANT: EPCS_TYPE STRING "EPCS64"
-- Retrieval info: CONSTANT: FLASH_RSTPIN STRING "FALSE"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
-- Retrieval info: CONSTANT: LPM_HINT STRING "UNUSED"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "altasmi_parallel"
-- Retrieval info: CONSTANT: PAGE_SIZE NUMERIC "1"
-- Retrieval info: CONSTANT: PORT_BULK_ERASE STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_DIE_ERASE STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_EN4B_ADDR STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_EX4B_ADDR STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_FAST_READ STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_ILLEGAL_ERASE STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_ILLEGAL_WRITE STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_RDID_OUT STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_READ_ADDRESS STRING "PORT_USED"
-- Retrieval info: CONSTANT: PORT_READ_DUMMYCLK STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_READ_RDID STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_READ_SID STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_READ_STATUS STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_SECTOR_ERASE STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_SECTOR_PROTECT STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_SHIFT_BYTES STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_WREN STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_WRITE STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: USE_ASMIBLOCK STRING "ON"
-- Retrieval info: CONSTANT: USE_EAB STRING "ON"
-- Retrieval info: CONSTANT: WRITE_DUMMY_CLK NUMERIC "0"
-- Retrieval info: USED_PORT: addr 0 0 24 0 INPUT NODEFVAL "addr[23..0]"
-- Retrieval info: CONNECT: @addr 0 0 24 0 addr 0 0 24 0
-- Retrieval info: USED_PORT: busy 0 0 0 0 OUTPUT NODEFVAL "busy"
-- Retrieval info: CONNECT: busy 0 0 0 0 @busy 0 0 0 0
-- Retrieval info: USED_PORT: clkin 0 0 0 0 INPUT NODEFVAL "clkin"
-- Retrieval info: CONNECT: @clkin 0 0 0 0 clkin 0 0 0 0
-- Retrieval info: USED_PORT: data_valid 0 0 0 0 OUTPUT NODEFVAL "data_valid"
-- Retrieval info: CONNECT: data_valid 0 0 0 0 @data_valid 0 0 0 0
-- Retrieval info: USED_PORT: dataout 0 0 8 0 OUTPUT NODEFVAL "dataout[7..0]"
-- Retrieval info: CONNECT: dataout 0 0 8 0 @dataout 0 0 8 0
-- Retrieval info: USED_PORT: rden 0 0 0 0 INPUT NODEFVAL "rden"
-- Retrieval info: CONNECT: @rden 0 0 0 0 rden 0 0 0 0
-- Retrieval info: USED_PORT: read 0 0 0 0 INPUT NODEFVAL "read"
-- Retrieval info: CONNECT: @read 0 0 0 0 read 0 0 0 0
-- Retrieval info: USED_PORT: read_address 0 0 24 0 OUTPUT NODEFVAL "read_address[23..0]"
-- Retrieval info: CONNECT: read_address 0 0 24 0 @read_address 0 0 24 0
-- Retrieval info: USED_PORT: reset 0 0 0 0 INPUT NODEFVAL "reset"
-- Retrieval info: CONNECT: @reset 0 0 0 0 reset 0 0 0 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL asmicont.vhd TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL asmicont.qip TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL asmicont.bsf TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL asmicont_inst.vhd TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL asmicont.inc TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL asmicont.cmp TRUE TRUE

-- megafunction wizard: %ALTASMI_PARALLEL%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: ALTASMI_PARALLEL 

-- ============================================================
-- File Name: asmicont.vhd
-- Megafunction Name(s):
-- 			ALTASMI_PARALLEL
--
-- Simulation Library Files(s):
-- 			
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 13.1.0 Build 162 10/23/2013 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2013 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


--altasmi_parallel CBX_AUTO_BLACKBOX="ALL" DATA_WIDTH="STANDARD" DEVICE_FAMILY="Cyclone V" EPCS_TYPE="EPCS64" PAGE_SIZE=1 PORT_BULK_ERASE="PORT_UNUSED" PORT_DIE_ERASE="PORT_UNUSED" PORT_EN4B_ADDR="PORT_UNUSED" PORT_EX4B_ADDR="PORT_UNUSED" PORT_FAST_READ="PORT_UNUSED" PORT_ILLEGAL_ERASE="PORT_UNUSED" PORT_ILLEGAL_WRITE="PORT_UNUSED" PORT_RDID_OUT="PORT_UNUSED" PORT_READ_ADDRESS="PORT_USED" PORT_READ_DUMMYCLK="PORT_UNUSED" PORT_READ_RDID="PORT_UNUSED" PORT_READ_SID="PORT_UNUSED" PORT_READ_STATUS="PORT_UNUSED" PORT_SECTOR_ERASE="PORT_UNUSED" PORT_SECTOR_PROTECT="PORT_UNUSED" PORT_SHIFT_BYTES="PORT_UNUSED" PORT_WREN="PORT_UNUSED" PORT_WRITE="PORT_UNUSED" USE_ASMIBLOCK="ON" USE_EAB="ON" WRITE_DUMMY_CLK=0 addr busy clkin data_valid dataout rden read read_address reset INTENDED_DEVICE_FAMILY="Cyclone V" ALTERA_INTERNAL_OPTIONS=SUPPRESS_DA_RULE_INTERNAL=C106
--VERSION_BEGIN 13.1 cbx_a_gray2bin 2013:10:23:18:05:48:SJ cbx_a_graycounter 2013:10:23:18:05:48:SJ cbx_altasmi_parallel 2013:10:23:18:05:48:SJ cbx_altdpram 2013:10:23:18:05:48:SJ cbx_altsyncram 2013:10:23:18:05:48:SJ cbx_arriav 2013:10:23:18:05:48:SJ cbx_cyclone 2013:10:23:18:05:48:SJ cbx_cycloneii 2013:10:23:18:05:48:SJ cbx_fifo_common 2013:10:23:18:05:48:SJ cbx_lpm_add_sub 2013:10:23:18:05:48:SJ cbx_lpm_compare 2013:10:23:18:05:48:SJ cbx_lpm_counter 2013:10:23:18:05:48:SJ cbx_lpm_decode 2013:10:23:18:05:48:SJ cbx_lpm_mux 2013:10:23:18:05:48:SJ cbx_mgl 2013:10:23:18:06:54:SJ cbx_nightfury 2013:10:23:18:05:48:SJ cbx_scfifo 2013:10:23:18:05:48:SJ cbx_stratix 2013:10:23:18:05:48:SJ cbx_stratixii 2013:10:23:18:05:48:SJ cbx_stratixiii 2013:10:23:18:05:48:SJ cbx_stratixv 2013:10:23:18:05:48:SJ cbx_util_mgl 2013:10:23:18:05:48:SJ  VERSION_END

 LIBRARY altera_mf;
 USE altera_mf.all;

 LIBRARY cyclonev;
 USE cyclonev.all;

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = a_graycounter 3 cyclonev_asmiblock 1 lpm_counter 1 lut 6 mux21 1 reg 91 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  asmicont_altasmi_parallel_qth2 IS 
	 PORT 
	 ( 
		 addr	:	IN  STD_LOGIC_VECTOR (23 DOWNTO 0);
		 busy	:	OUT  STD_LOGIC;
		 clkin	:	IN  STD_LOGIC;
		 data_valid	:	OUT  STD_LOGIC;
		 dataout	:	OUT  STD_LOGIC_VECTOR (7 DOWNTO 0);
		 rden	:	IN  STD_LOGIC;
		 read	:	IN  STD_LOGIC := '0';
		 read_address	:	OUT  STD_LOGIC_VECTOR (23 DOWNTO 0);
		 reset	:	IN  STD_LOGIC := '0'
	 ); 
 END asmicont_altasmi_parallel_qth2;

 ARCHITECTURE RTL OF asmicont_altasmi_parallel_qth2 IS

	 ATTRIBUTE synthesis_clearbox : natural;
	 ATTRIBUTE synthesis_clearbox OF RTL : ARCHITECTURE IS 2;
	 ATTRIBUTE ALTERA_ATTRIBUTE : string;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF RTL : ARCHITECTURE IS "SUPPRESS_DA_RULE_INTERNAL=C106";

	 SIGNAL  wire_addbyte_cntr_w_lg_w_q_range144w149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addbyte_cntr_w_lg_w_q_range147w148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addbyte_cntr_clk_en	:	STD_LOGIC;
	 SIGNAL  wire_stage_cntr_w143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addbyte_cntr_clock	:	STD_LOGIC;
	 SIGNAL  wire_addbyte_cntr_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_addbyte_cntr_sclr	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_end_operation86w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addbyte_cntr_w_q_range147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addbyte_cntr_w_q_range144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_gen_cntr_w_lg_w_q_range99w100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_gen_cntr_w_lg_w_q_range97w98w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_gen_cntr_clk_en	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_w_lg_in_operation26w27w28w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_gen_cntr_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_gen_cntr_sclr	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_end1_cyc_reg_in_wire29w30w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_gen_cntr_w_q_range97w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_gen_cntr_w_q_range99w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w325w326w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w325w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w330w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range89w92w322w323w324w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range89w92w327w328w329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range89w90w91w336w337w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range89w94w413w414w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range89w92w322w323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range89w92w347w348w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range89w92w327w328w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range89w90w91w336w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range89w94w413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range89w92w322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range89w92w347w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range89w92w327w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range89w92w140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range89w92w320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range88w93w119w120w121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range88w93w119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range89w90w91w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_q_range89w94w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_q_range89w92w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range88w93w119w120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_q_range88w93w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_q_range89w90w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_clk_en	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_w_lg_w82w83w84w85w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_sclr	:	STD_LOGIC;
	 SIGNAL  wire_stage_cntr_w_q_range88w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_q_range89w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_arriav_asmiblock2_data1in	:	STD_LOGIC;
	 SIGNAL  wire_vcc	:	STD_LOGIC;
	 SIGNAL	 add_msb_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_add_msb_reg_ena	:	STD_LOGIC;
	 SIGNAL	 add_rollover_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_addr_reg_d	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL	 addr_reg	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_addr_reg_ena	:	STD_LOGIC_VECTOR(23 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_q_range386w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL	 wire_asmi_opcode_reg_d	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL	 asmi_opcode_reg	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_asmi_opcode_reg_ena	:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	 SIGNAL  wire_asmi_opcode_reg_w_q_range154w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL	 busy_det_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 clr_read_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 clr_read_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dvalid_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_dvalid_reg_ena	:	STD_LOGIC;
	 SIGNAL	 wire_dvalid_reg_sclr	:	STD_LOGIC;
	 SIGNAL	 dvalid_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 end1_cyc_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 end1_cyc_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 end_op_hdlyreg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 end_op_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 end_rbyte_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_end_rbyte_reg_ena	:	STD_LOGIC;
	 SIGNAL	 wire_end_rbyte_reg_sclr	:	STD_LOGIC;
	 SIGNAL	 end_read_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 ncs_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_ncs_reg_sclr	:	STD_LOGIC;
	 SIGNAL  wire_ncs_reg_w_lg_q373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 wire_read_add_reg_d	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL	 read_add_reg	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_read_add_reg_ena	:	STD_LOGIC_VECTOR(23 DOWNTO 0);
	 SIGNAL	 wire_read_data_reg_d	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL	 read_data_reg	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_read_data_reg_ena	:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	 SIGNAL	 wire_read_dout_reg_d	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL	 read_dout_reg	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_read_dout_reg_ena	:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	 SIGNAL	 read_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_read_reg_ena	:	STD_LOGIC;
	 SIGNAL	 shift_op_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 stage2_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 stage3_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 stage4_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_read_add_cntr_clk_en	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_w_lg_rden_wire476w477w478w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_read_add_cntr_data	:	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  wire_read_add_cntr_q	:	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  wire_read_add_cntr_sload	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_rden_wire476w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	wire_mux211_dataout	:	STD_LOGIC;
	 SIGNAL  wire_w273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w213w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w271w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w206w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w470w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode170w171w172w257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode170w171w172w173w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode175w176w177w259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode175w176w177w178w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode209w210w211w212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode180w181w182w261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode180w181w182w183w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode221w222w223w279w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode221w222w223w224w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode202w203w204w205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_read352w353w354w355w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_read400w467w468w469w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_sec_erase40w409w410w411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode170w171w172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode175w176w177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode185w190w265w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode185w190w191w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode185w186w263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode185w186w187w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode209w210w211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode180w181w182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode221w222w223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode202w203w204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_read352w353w354w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_read352w353w412w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_read400w467w468w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_sec_erase40w409w410w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_4baddr162w163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_ex4baddr157w158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read_stat109w110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_write193w194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_write49w331w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_end_read_byte474w486w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode164w253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode164w165w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode159w251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode159w160w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode195w267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode195w196w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode170w171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode175w176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode215w275w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode215w216w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode218w277w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode218w219w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode198w269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode198w199w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode226w281w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode226w227w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode229w283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode229w230w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode185w190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode185w186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode209w210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode180w181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode221w222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode167w255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode167w168w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode202w203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_stage3_wire31w32w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_start_poll338w339w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read352w353w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_write58w102w103w116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_write58w59w401w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read400w467w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read_rdid111w112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_sec_erase40w409w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_rden_wire405w406w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_addr_overdie395w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_addr_overdie385w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_4baddr162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_bulk_erase332w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_ex4baddr157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read_nonvolatile318w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read_stat109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_write193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_write56w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_write49w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_read_byte474w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode215w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode229w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_not_busy397w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_not_busy389w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_opcode155w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage3_wire403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage3_wire434w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage3_wire41w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage3_wire31w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage3_wire387w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage4_wire436w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage4_wire404w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_start_poll338w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_write49w350w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w105w106w107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_addr_overdie499w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_busy_wire1w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_clkin_wire87w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_fast_read351w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_memadd418w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_polling189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read352w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read_rdid37w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read_stat38w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read_volatile201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_wren39w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_write_volatile208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_add_cycle69w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_fast_read63w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_operation485w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_ophdly25w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_pgwr_data48w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_read66w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rden_wire501w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_rdid_wire7w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_sid_wire6w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_sec_protect_wire5w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_st_busy_wire113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_start_poll108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_pagewr_buf_not_empty_range54w55w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode229w283w284w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode229w230w231w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_write58w59w401w402w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_rden_wire405w406w407w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_not_busy397w398w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_not_busy389w390w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_stage4_wire436w437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode229w283w284w285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode229w230w231w232w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_rden_wire405w406w407w408w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_not_busy389w390w391w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w233w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w286w287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w233w234w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w286w287w288w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w233w234w235w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w286w287w288w289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w233w234w235w236w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w286w287w288w289w290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w233w234w235w236w237w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w286w287w288w289w290w291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w233w234w235w236w237w238w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w239w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w292w293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w239w240w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w292w293w294w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w239w240w241w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w292w293w294w295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w239w240w241w242w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w292w293w294w295w296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w239w240w241w242w243w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w292w293w294w295w296w297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w239w240w241w242w243w244w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w245w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w298w299w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w245w246w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w245w246w247w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w137w138w139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w137w138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w105w106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_read400w421w422w423w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_read_sid133w134w135w136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_write58w102w103w104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_read400w421w422w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_read_sid133w134w135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_read_stat431w432w433w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_write58w102w103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read400w435w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read400w421w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read_sid133w134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read_stat431w432w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_write58w102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_write58w59w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_data0out_wire439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_4baddr334w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_ex4baddr333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read400w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read_rdid111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read_sid133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read_stat431w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_sec_erase40w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_wren335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_write58w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rden_wire405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  add_rollover :	STD_LOGIC;
	 SIGNAL  addr_overdie :	STD_LOGIC;
	 SIGNAL  addr_overdie_pos :	STD_LOGIC;
	 SIGNAL  addr_reg_overdie :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  b4addr_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  berase_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  busy_wire :	STD_LOGIC;
	 SIGNAL  clkin_wire :	STD_LOGIC;
	 SIGNAL  clr_addmsb_wire :	STD_LOGIC;
	 SIGNAL  clr_endrbyte_wire :	STD_LOGIC;
	 SIGNAL  clr_read_wire :	STD_LOGIC;
	 SIGNAL  clr_read_wire2 :	STD_LOGIC;
	 SIGNAL  clr_write_wire2 :	STD_LOGIC;
	 SIGNAL  data0out_wire :	STD_LOGIC;
	 SIGNAL  data_valid_wire :	STD_LOGIC;
	 SIGNAL  dataoe_wire :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  dataout_wire :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  derase_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  do_4baddr :	STD_LOGIC;
	 SIGNAL  do_bulk_erase :	STD_LOGIC;
	 SIGNAL  do_die_erase :	STD_LOGIC;
	 SIGNAL  do_ex4baddr :	STD_LOGIC;
	 SIGNAL  do_fast_read :	STD_LOGIC;
	 SIGNAL  do_fread_epcq :	STD_LOGIC;
	 SIGNAL  do_freadwrv_polling :	STD_LOGIC;
	 SIGNAL  do_memadd :	STD_LOGIC;
	 SIGNAL  do_polling :	STD_LOGIC;
	 SIGNAL  do_read :	STD_LOGIC;
	 SIGNAL  do_read_nonvolatile :	STD_LOGIC;
	 SIGNAL  do_read_rdid :	STD_LOGIC;
	 SIGNAL  do_read_sid :	STD_LOGIC;
	 SIGNAL  do_read_stat :	STD_LOGIC;
	 SIGNAL  do_read_volatile :	STD_LOGIC;
	 SIGNAL  do_sec_erase :	STD_LOGIC;
	 SIGNAL  do_sec_prot :	STD_LOGIC;
	 SIGNAL  do_sprot_polling :	STD_LOGIC;
	 SIGNAL  do_wait_dummyclk :	STD_LOGIC;
	 SIGNAL  do_wren :	STD_LOGIC;
	 SIGNAL  do_write :	STD_LOGIC;
	 SIGNAL  do_write_polling :	STD_LOGIC;
	 SIGNAL  do_write_volatile :	STD_LOGIC;
	 SIGNAL  end1_cyc_gen_cntr_wire :	STD_LOGIC;
	 SIGNAL  end1_cyc_normal_in_wire :	STD_LOGIC;
	 SIGNAL  end1_cyc_reg_in_wire :	STD_LOGIC;
	 SIGNAL  end_add_cycle :	STD_LOGIC;
	 SIGNAL  end_add_cycle_mux_datab_wire :	STD_LOGIC;
	 SIGNAL  end_fast_read :	STD_LOGIC;
	 SIGNAL  end_one_cyc_pos :	STD_LOGIC;
	 SIGNAL  end_one_cycle :	STD_LOGIC;
	 SIGNAL  end_op_wire :	STD_LOGIC;
	 SIGNAL  end_operation :	STD_LOGIC;
	 SIGNAL  end_ophdly :	STD_LOGIC;
	 SIGNAL  end_pgwr_data :	STD_LOGIC;
	 SIGNAL  end_read :	STD_LOGIC;
	 SIGNAL  end_read_byte :	STD_LOGIC;
	 SIGNAL  exb4addr_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  fast_read_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  freadwrv_sdoin :	STD_LOGIC;
	 SIGNAL  in_operation :	STD_LOGIC;
	 SIGNAL  load_opcode :	STD_LOGIC;
	 SIGNAL  memadd_sdoin :	STD_LOGIC;
	 SIGNAL  ncs_reg_ena_wire :	STD_LOGIC;
	 SIGNAL  not_busy :	STD_LOGIC;
	 SIGNAL  oe_wire :	STD_LOGIC;
	 SIGNAL  pagewr_buf_not_empty :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  rden_wire :	STD_LOGIC;
	 SIGNAL  rdid_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  rdummyclk_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  read_data_reg_in_wire :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  read_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  read_rdid_wire :	STD_LOGIC;
	 SIGNAL  read_sid_wire :	STD_LOGIC;
	 SIGNAL  read_wire :	STD_LOGIC;
	 SIGNAL  rflagstat_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  rnvdummyclk_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  rsid_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  rsid_sdoin :	STD_LOGIC;
	 SIGNAL  rstat_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  scein_wire :	STD_LOGIC;
	 SIGNAL  sdoin_wire :	STD_LOGIC;
	 SIGNAL  sec_protect_wire :	STD_LOGIC;
	 SIGNAL  secprot_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  secprot_sdoin :	STD_LOGIC;
	 SIGNAL  serase_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  shift_opcode :	STD_LOGIC;
	 SIGNAL  shift_opdata :	STD_LOGIC;
	 SIGNAL  shift_pgwr_data :	STD_LOGIC;
	 SIGNAL  st_busy_wire :	STD_LOGIC;
	 SIGNAL  stage2_wire :	STD_LOGIC;
	 SIGNAL  stage3_wire :	STD_LOGIC;
	 SIGNAL  stage4_wire :	STD_LOGIC;
	 SIGNAL  start_frpoll :	STD_LOGIC;
	 SIGNAL  start_poll :	STD_LOGIC;
	 SIGNAL  start_sppoll :	STD_LOGIC;
	 SIGNAL  start_wrpoll :	STD_LOGIC;
	 SIGNAL  to_sdoin_wire :	STD_LOGIC;
	 SIGNAL  wren_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wren_wire :	STD_LOGIC;
	 SIGNAL  write_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  write_prot_true :	STD_LOGIC;
	 SIGNAL  write_sdoin :	STD_LOGIC;
	 SIGNAL  wrvolatile_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_addr_range396w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_addr_range388w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_addr_reg_overdie_range394w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_addr_reg_overdie_range384w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_b4addr_opcode_range252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_b4addr_opcode_range161w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_berase_opcode_range256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_berase_opcode_range169w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_dataout_wire_range438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_derase_opcode_range258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_derase_opcode_range174w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_exb4addr_opcode_range250w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exb4addr_opcode_range156w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_fast_read_opcode_range274w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_fast_read_opcode_range214w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_pagewr_buf_not_empty_range54w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rdid_opcode_range280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rdid_opcode_range225w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_rdummyclk_opcode_range272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rdummyclk_opcode_range207w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_read_opcode_range276w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_read_opcode_range217w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_rflagstat_opcode_range262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rflagstat_opcode_range184w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_rnvdummyclk_opcode_range268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rnvdummyclk_opcode_range197w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_rsid_opcode_range282w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rsid_opcode_range228w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_rstat_opcode_range264w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rstat_opcode_range188w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_secprot_opcode_range278w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_secprot_opcode_range220w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_serase_opcode_range260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_serase_opcode_range179w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_wren_opcode_range254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_wren_opcode_range166w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_write_opcode_range266w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_write_opcode_range192w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_wrvolatile_opcode_range270w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_wrvolatile_opcode_range200w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 COMPONENT  a_graycounter
	 GENERIC 
	 (
		PVALUE	:	NATURAL := 0;
		WIDTH	:	NATURAL := 8;
		lpm_type	:	STRING := "a_graycounter"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clk_en	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC;
		cnt_en	:	IN STD_LOGIC := '1';
		q	:	OUT STD_LOGIC_VECTOR(width-1 DOWNTO 0);
		qbin	:	OUT STD_LOGIC_VECTOR(width-1 DOWNTO 0);
		sclr	:	IN STD_LOGIC := '0';
		updown	:	IN STD_LOGIC := '1'
	 ); 
	 END COMPONENT;
	 COMPONENT  cyclonev_asmiblock
	 PORT
	 ( 
		data0in	:	OUT STD_LOGIC;
		data0oe	:	IN STD_LOGIC := '0';
		data0out	:	IN STD_LOGIC := '0';
		data1in	:	OUT STD_LOGIC;
		data1oe	:	IN STD_LOGIC := '0';
		data1out	:	IN STD_LOGIC := '0';
		data2in	:	OUT STD_LOGIC;
		data2oe	:	IN STD_LOGIC := '0';
		data2out	:	IN STD_LOGIC := '0';
		data3in	:	OUT STD_LOGIC;
		data3oe	:	IN STD_LOGIC := '0';
		data3out	:	IN STD_LOGIC := '0';
		dclk	:	IN STD_LOGIC;
		oe	:	IN STD_LOGIC := '0';
		sce	:	IN STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_counter
	 GENERIC 
	 (
		lpm_avalue	:	STRING := "0";
		lpm_direction	:	STRING := "DEFAULT";
		lpm_modulus	:	NATURAL := 0;
		lpm_port_updown	:	STRING := "PORT_CONNECTIVITY";
		lpm_pvalue	:	STRING := "0";
		lpm_svalue	:	STRING := "0";
		lpm_width	:	NATURAL;
		lpm_type	:	STRING := "lpm_counter"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aload	:	IN STD_LOGIC := '0';
		aset	:	IN STD_LOGIC := '0';
		cin	:	IN STD_LOGIC := '1';
		clk_en	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC;
		cnt_en	:	IN STD_LOGIC := '1';
		cout	:	OUT STD_LOGIC;
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		eq	:	OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		sclr	:	IN STD_LOGIC := '0';
		sload	:	IN STD_LOGIC := '0';
		sset	:	IN STD_LOGIC := '0';
		updown	:	IN STD_LOGIC := '1'
	 ); 
	 END COMPONENT;
 BEGIN

	wire_vcc <= '1';
	wire_w273w(0) <= wire_w_lg_w_lg_w_lg_w_lg_load_opcode209w210w211w212w(0) AND wire_w_rdummyclk_opcode_range272w(0);
	loop0 : FOR i IN 0 TO 6 GENERATE 
		wire_w213w(i) <= wire_w_lg_w_lg_w_lg_w_lg_load_opcode209w210w211w212w(0) AND wire_w_rdummyclk_opcode_range207w(i);
	END GENERATE loop0;
	wire_w271w(0) <= wire_w_lg_w_lg_w_lg_w_lg_load_opcode202w203w204w205w(0) AND wire_w_wrvolatile_opcode_range270w(0);
	loop1 : FOR i IN 0 TO 6 GENERATE 
		wire_w206w(i) <= wire_w_lg_w_lg_w_lg_w_lg_load_opcode202w203w204w205w(0) AND wire_w_wrvolatile_opcode_range200w(i);
	END GENERATE loop1;
	wire_w470w(0) <= wire_w_lg_w_lg_w_lg_w_lg_do_read400w467w468w469w(0) AND end_read_byte;
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode170w171w172w257w(0) <= wire_w_lg_w_lg_w_lg_load_opcode170w171w172w(0) AND wire_w_berase_opcode_range256w(0);
	loop2 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_load_opcode170w171w172w173w(i) <= wire_w_lg_w_lg_w_lg_load_opcode170w171w172w(0) AND wire_w_berase_opcode_range169w(i);
	END GENERATE loop2;
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode175w176w177w259w(0) <= wire_w_lg_w_lg_w_lg_load_opcode175w176w177w(0) AND wire_w_derase_opcode_range258w(0);
	loop3 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_load_opcode175w176w177w178w(i) <= wire_w_lg_w_lg_w_lg_load_opcode175w176w177w(0) AND wire_w_derase_opcode_range174w(i);
	END GENERATE loop3;
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode209w210w211w212w(0) <= wire_w_lg_w_lg_w_lg_load_opcode209w210w211w(0) AND wire_w_lg_do_read_stat38w(0);
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode180w181w182w261w(0) <= wire_w_lg_w_lg_w_lg_load_opcode180w181w182w(0) AND wire_w_serase_opcode_range260w(0);
	loop4 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_load_opcode180w181w182w183w(i) <= wire_w_lg_w_lg_w_lg_load_opcode180w181w182w(0) AND wire_w_serase_opcode_range179w(i);
	END GENERATE loop4;
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode221w222w223w279w(0) <= wire_w_lg_w_lg_w_lg_load_opcode221w222w223w(0) AND wire_w_secprot_opcode_range278w(0);
	loop5 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_load_opcode221w222w223w224w(i) <= wire_w_lg_w_lg_w_lg_load_opcode221w222w223w(0) AND wire_w_secprot_opcode_range220w(i);
	END GENERATE loop5;
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode202w203w204w205w(0) <= wire_w_lg_w_lg_w_lg_load_opcode202w203w204w(0) AND wire_w_lg_do_read_stat38w(0);
	wire_w_lg_w_lg_w_lg_w_lg_do_read352w353w354w355w(0) <= wire_w_lg_w_lg_w_lg_do_read352w353w354w(0) AND end_one_cycle;
	wire_w_lg_w_lg_w_lg_w_lg_do_read400w467w468w469w(0) <= wire_w_lg_w_lg_w_lg_do_read400w467w468w(0) AND end_one_cyc_pos;
	wire_w_lg_w_lg_w_lg_w_lg_do_sec_erase40w409w410w411w(0) <= wire_w_lg_w_lg_w_lg_do_sec_erase40w409w410w(0) AND end_operation;
	wire_w_lg_w_lg_w_lg_load_opcode170w171w172w(0) <= wire_w_lg_w_lg_load_opcode170w171w(0) AND wire_w_lg_do_read_stat38w(0);
	wire_w_lg_w_lg_w_lg_load_opcode175w176w177w(0) <= wire_w_lg_w_lg_load_opcode175w176w(0) AND wire_w_lg_do_read_stat38w(0);
	wire_w_lg_w_lg_w_lg_load_opcode185w190w265w(0) <= wire_w_lg_w_lg_load_opcode185w190w(0) AND wire_w_rstat_opcode_range264w(0);
	loop6 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_load_opcode185w190w191w(i) <= wire_w_lg_w_lg_load_opcode185w190w(0) AND wire_w_rstat_opcode_range188w(i);
	END GENERATE loop6;
	wire_w_lg_w_lg_w_lg_load_opcode185w186w263w(0) <= wire_w_lg_w_lg_load_opcode185w186w(0) AND wire_w_rflagstat_opcode_range262w(0);
	loop7 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_load_opcode185w186w187w(i) <= wire_w_lg_w_lg_load_opcode185w186w(0) AND wire_w_rflagstat_opcode_range184w(i);
	END GENERATE loop7;
	wire_w_lg_w_lg_w_lg_load_opcode209w210w211w(0) <= wire_w_lg_w_lg_load_opcode209w210w(0) AND wire_w_lg_do_wren39w(0);
	wire_w_lg_w_lg_w_lg_load_opcode180w181w182w(0) <= wire_w_lg_w_lg_load_opcode180w181w(0) AND wire_w_lg_do_read_stat38w(0);
	wire_w_lg_w_lg_w_lg_load_opcode221w222w223w(0) <= wire_w_lg_w_lg_load_opcode221w222w(0) AND wire_w_lg_do_read_stat38w(0);
	wire_w_lg_w_lg_w_lg_load_opcode202w203w204w(0) <= wire_w_lg_w_lg_load_opcode202w203w(0) AND wire_w_lg_do_wren39w(0);
	wire_w_lg_w_lg_w_lg_do_read352w353w354w(0) <= wire_w_lg_w_lg_do_read352w353w(0) AND wire_w_lg_w_lg_do_write49w350w(0);
	wire_w_lg_w_lg_w_lg_do_read352w353w412w(0) <= wire_w_lg_w_lg_do_read352w353w(0) AND clr_write_wire2;
	wire_w_lg_w_lg_w_lg_do_read400w467w468w(0) <= wire_w_lg_w_lg_do_read400w467w(0) AND wire_stage_cntr_w_lg_w_q_range88w93w(0);
	wire_w_lg_w_lg_w_lg_do_sec_erase40w409w410w(0) <= wire_w_lg_w_lg_do_sec_erase40w409w(0) AND wire_w_lg_do_read_stat38w(0);
	wire_w_lg_w_lg_do_4baddr162w163w(0) <= wire_w_lg_do_4baddr162w(0) AND wire_w_lg_do_wren39w(0);
	wire_w_lg_w_lg_do_ex4baddr157w158w(0) <= wire_w_lg_do_ex4baddr157w(0) AND wire_w_lg_do_wren39w(0);
	wire_w_lg_w_lg_do_read_stat109w110w(0) <= wire_w_lg_do_read_stat109w(0) AND wire_w_lg_w_lg_w105w106w107w(0);
	wire_w_lg_w_lg_do_write193w194w(0) <= wire_w_lg_do_write193w(0) AND wire_w_lg_do_wren39w(0);
	wire_w_lg_w_lg_do_write49w331w(0) <= wire_w_lg_do_write49w(0) AND end_pgwr_data;
	wire_w_lg_w_lg_end_read_byte474w486w(0) <= wire_w_lg_end_read_byte474w(0) AND wire_w_lg_end_operation485w(0);
	wire_w_lg_w_lg_load_opcode164w253w(0) <= wire_w_lg_load_opcode164w(0) AND wire_w_b4addr_opcode_range252w(0);
	loop8 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode164w165w(i) <= wire_w_lg_load_opcode164w(0) AND wire_w_b4addr_opcode_range161w(i);
	END GENERATE loop8;
	wire_w_lg_w_lg_load_opcode159w251w(0) <= wire_w_lg_load_opcode159w(0) AND wire_w_exb4addr_opcode_range250w(0);
	loop9 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode159w160w(i) <= wire_w_lg_load_opcode159w(0) AND wire_w_exb4addr_opcode_range156w(i);
	END GENERATE loop9;
	wire_w_lg_w_lg_load_opcode195w267w(0) <= wire_w_lg_load_opcode195w(0) AND wire_w_write_opcode_range266w(0);
	loop10 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode195w196w(i) <= wire_w_lg_load_opcode195w(0) AND wire_w_write_opcode_range192w(i);
	END GENERATE loop10;
	wire_w_lg_w_lg_load_opcode170w171w(0) <= wire_w_lg_load_opcode170w(0) AND wire_w_lg_do_wren39w(0);
	wire_w_lg_w_lg_load_opcode175w176w(0) <= wire_w_lg_load_opcode175w(0) AND wire_w_lg_do_wren39w(0);
	wire_w_lg_w_lg_load_opcode215w275w(0) <= wire_w_lg_load_opcode215w(0) AND wire_w_fast_read_opcode_range274w(0);
	loop11 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode215w216w(i) <= wire_w_lg_load_opcode215w(0) AND wire_w_fast_read_opcode_range214w(i);
	END GENERATE loop11;
	wire_w_lg_w_lg_load_opcode218w277w(0) <= wire_w_lg_load_opcode218w(0) AND wire_w_read_opcode_range276w(0);
	loop12 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode218w219w(i) <= wire_w_lg_load_opcode218w(0) AND wire_w_read_opcode_range217w(i);
	END GENERATE loop12;
	wire_w_lg_w_lg_load_opcode198w269w(0) <= wire_w_lg_load_opcode198w(0) AND wire_w_rnvdummyclk_opcode_range268w(0);
	loop13 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode198w199w(i) <= wire_w_lg_load_opcode198w(0) AND wire_w_rnvdummyclk_opcode_range197w(i);
	END GENERATE loop13;
	wire_w_lg_w_lg_load_opcode226w281w(0) <= wire_w_lg_load_opcode226w(0) AND wire_w_rdid_opcode_range280w(0);
	loop14 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode226w227w(i) <= wire_w_lg_load_opcode226w(0) AND wire_w_rdid_opcode_range225w(i);
	END GENERATE loop14;
	wire_w_lg_w_lg_load_opcode229w283w(0) <= wire_w_lg_load_opcode229w(0) AND wire_w_rsid_opcode_range282w(0);
	loop15 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode229w230w(i) <= wire_w_lg_load_opcode229w(0) AND wire_w_rsid_opcode_range228w(i);
	END GENERATE loop15;
	wire_w_lg_w_lg_load_opcode185w190w(0) <= wire_w_lg_load_opcode185w(0) AND wire_w_lg_do_polling189w(0);
	wire_w_lg_w_lg_load_opcode185w186w(0) <= wire_w_lg_load_opcode185w(0) AND do_polling;
	wire_w_lg_w_lg_load_opcode209w210w(0) <= wire_w_lg_load_opcode209w(0) AND wire_w_lg_do_write_volatile208w(0);
	wire_w_lg_w_lg_load_opcode180w181w(0) <= wire_w_lg_load_opcode180w(0) AND wire_w_lg_do_wren39w(0);
	wire_w_lg_w_lg_load_opcode221w222w(0) <= wire_w_lg_load_opcode221w(0) AND wire_w_lg_do_wren39w(0);
	wire_w_lg_w_lg_load_opcode167w255w(0) <= wire_w_lg_load_opcode167w(0) AND wire_w_wren_opcode_range254w(0);
	loop16 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode167w168w(i) <= wire_w_lg_load_opcode167w(0) AND wire_w_wren_opcode_range166w(i);
	END GENERATE loop16;
	wire_w_lg_w_lg_load_opcode202w203w(0) <= wire_w_lg_load_opcode202w(0) AND wire_w_lg_do_read_volatile201w(0);
	wire_w_lg_w_lg_stage3_wire31w32w(0) <= wire_w_lg_stage3_wire31w(0) AND do_wait_dummyclk;
	wire_w_lg_w_lg_start_poll338w339w(0) <= wire_w_lg_start_poll338w(0) AND do_polling;
	wire_w_lg_w_lg_do_read352w353w(0) <= wire_w_lg_do_read352w(0) AND wire_w_lg_do_fast_read351w(0);
	wire_w_lg_w_lg_w_lg_w_lg_do_write58w102w103w116w(0) <= wire_w_lg_w_lg_w_lg_do_write58w102w103w(0) AND write_prot_true;
	wire_w_lg_w_lg_w_lg_do_write58w59w401w(0) <= wire_w_lg_w_lg_do_write58w59w(0) AND do_memadd;
	wire_w_lg_w_lg_do_read400w467w(0) <= wire_w_lg_do_read400w(0) AND wire_stage_cntr_w_q_range89w(0);
	wire_w_lg_w_lg_do_read_rdid111w112w(0) <= wire_w_lg_do_read_rdid111w(0) AND end_op_wire;
	wire_w_lg_w_lg_do_sec_erase40w409w(0) <= wire_w_lg_do_sec_erase40w(0) AND wire_w_lg_do_wren39w(0);
	wire_w_lg_w_lg_rden_wire405w406w(0) <= wire_w_lg_rden_wire405w(0) AND not_busy;
	wire_w_lg_addr_overdie395w(0) <= addr_overdie AND wire_w_addr_reg_overdie_range394w(0);
	loop17 : FOR i IN 0 TO 22 GENERATE 
		wire_w_lg_addr_overdie385w(i) <= addr_overdie AND wire_w_addr_reg_overdie_range384w(i);
	END GENERATE loop17;
	wire_w_lg_do_4baddr162w(0) <= do_4baddr AND wire_w_lg_do_read_stat38w(0);
	wire_w_lg_do_bulk_erase332w(0) <= do_bulk_erase AND wire_w_lg_do_read_stat38w(0);
	wire_w_lg_do_ex4baddr157w(0) <= do_ex4baddr AND wire_w_lg_do_read_stat38w(0);
	wire_w_lg_do_read_nonvolatile318w(0) <= do_read_nonvolatile AND wire_addbyte_cntr_w_q_range144w(0);
	wire_w_lg_do_read_stat109w(0) <= do_read_stat AND wire_w_lg_start_poll108w(0);
	wire_w_lg_do_write193w(0) <= do_write AND wire_w_lg_do_read_stat38w(0);
	wire_w_lg_do_write56w(0) <= do_write AND wire_w_lg_w_pagewr_buf_not_empty_range54w55w(0);
	wire_w_lg_do_write49w(0) <= do_write AND shift_pgwr_data;
	wire_w_lg_end_read_byte474w(0) <= end_read_byte AND end_one_cyc_pos;
	wire_w_lg_load_opcode164w(0) <= load_opcode AND wire_w_lg_w_lg_do_4baddr162w163w(0);
	wire_w_lg_load_opcode159w(0) <= load_opcode AND wire_w_lg_w_lg_do_ex4baddr157w158w(0);
	wire_w_lg_load_opcode195w(0) <= load_opcode AND wire_w_lg_w_lg_do_write193w194w(0);
	wire_w_lg_load_opcode170w(0) <= load_opcode AND do_bulk_erase;
	wire_w_lg_load_opcode175w(0) <= load_opcode AND do_die_erase;
	wire_w_lg_load_opcode215w(0) <= load_opcode AND do_fast_read;
	wire_w_lg_load_opcode218w(0) <= load_opcode AND do_read;
	wire_w_lg_load_opcode198w(0) <= load_opcode AND do_read_nonvolatile;
	wire_w_lg_load_opcode226w(0) <= load_opcode AND do_read_rdid;
	wire_w_lg_load_opcode229w(0) <= load_opcode AND do_read_sid;
	wire_w_lg_load_opcode185w(0) <= load_opcode AND do_read_stat;
	wire_w_lg_load_opcode209w(0) <= load_opcode AND do_read_volatile;
	wire_w_lg_load_opcode180w(0) <= load_opcode AND do_sec_erase;
	wire_w_lg_load_opcode221w(0) <= load_opcode AND do_sec_prot;
	wire_w_lg_load_opcode167w(0) <= load_opcode AND do_wren;
	wire_w_lg_load_opcode202w(0) <= load_opcode AND do_write_volatile;
	wire_w_lg_not_busy397w(0) <= not_busy AND wire_w_addr_range396w(0);
	loop18 : FOR i IN 0 TO 22 GENERATE 
		wire_w_lg_not_busy389w(i) <= not_busy AND wire_w_addr_range388w(i);
	END GENERATE loop18;
	loop19 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_shift_opcode155w(i) <= shift_opcode AND wire_asmi_opcode_reg_w_q_range154w(i);
	END GENERATE loop19;
	wire_w_lg_stage3_wire403w(0) <= stage3_wire AND wire_w_lg_w_lg_w_lg_w_lg_do_write58w59w401w402w(0);
	wire_w_lg_stage3_wire434w(0) <= stage3_wire AND wire_w_lg_w_lg_w_lg_do_read_stat431w432w433w(0);
	wire_w_lg_stage3_wire41w(0) <= stage3_wire AND wire_w_lg_do_sec_erase40w(0);
	wire_w_lg_stage3_wire31w(0) <= stage3_wire AND do_fast_read;
	loop20 : FOR i IN 0 TO 22 GENERATE 
		wire_w_lg_stage3_wire387w(i) <= stage3_wire AND wire_addr_reg_w_q_range386w(i);
	END GENERATE loop20;
	wire_w_lg_stage4_wire436w(0) <= stage4_wire AND wire_w_lg_w_lg_do_read400w435w(0);
	wire_w_lg_stage4_wire404w(0) <= stage4_wire AND addr_overdie;
	wire_w_lg_start_poll338w(0) <= start_poll AND do_read_stat;
	wire_w_lg_w_lg_do_write49w350w(0) <= NOT wire_w_lg_do_write49w(0);
	wire_w_lg_w_lg_w105w106w107w(0) <= NOT wire_w_lg_w105w106w(0);
	wire_w_lg_addr_overdie499w(0) <= NOT addr_overdie;
	wire_w_lg_busy_wire1w(0) <= NOT busy_wire;
	wire_w_lg_clkin_wire87w(0) <= NOT clkin_wire;
	wire_w_lg_do_fast_read351w(0) <= NOT do_fast_read;
	wire_w_lg_do_memadd418w(0) <= NOT do_memadd;
	wire_w_lg_do_polling189w(0) <= NOT do_polling;
	wire_w_lg_do_read352w(0) <= NOT do_read;
	wire_w_lg_do_read_rdid37w(0) <= NOT do_read_rdid;
	wire_w_lg_do_read_stat38w(0) <= NOT do_read_stat;
	wire_w_lg_do_read_volatile201w(0) <= NOT do_read_volatile;
	wire_w_lg_do_wren39w(0) <= NOT do_wren;
	wire_w_lg_do_write_volatile208w(0) <= NOT do_write_volatile;
	wire_w_lg_end_add_cycle69w(0) <= NOT end_add_cycle;
	wire_w_lg_end_fast_read63w(0) <= NOT end_fast_read;
	wire_w_lg_end_operation485w(0) <= NOT end_operation;
	wire_w_lg_end_ophdly25w(0) <= NOT end_ophdly;
	wire_w_lg_end_pgwr_data48w(0) <= NOT end_pgwr_data;
	wire_w_lg_end_read66w(0) <= NOT end_read;
	wire_w_lg_rden_wire501w(0) <= NOT rden_wire;
	wire_w_lg_read_rdid_wire7w(0) <= NOT read_rdid_wire;
	wire_w_lg_read_sid_wire6w(0) <= NOT read_sid_wire;
	wire_w_lg_sec_protect_wire5w(0) <= NOT sec_protect_wire;
	wire_w_lg_st_busy_wire113w(0) <= NOT st_busy_wire;
	wire_w_lg_start_poll108w(0) <= NOT start_poll;
	wire_w_lg_w_pagewr_buf_not_empty_range54w55w(0) <= NOT wire_w_pagewr_buf_not_empty_range54w(0);
	wire_w_lg_w_lg_w_lg_load_opcode229w283w284w(0) <= wire_w_lg_w_lg_load_opcode229w283w(0) OR wire_w_lg_w_lg_load_opcode226w281w(0);
	loop21 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_load_opcode229w230w231w(i) <= wire_w_lg_w_lg_load_opcode229w230w(i) OR wire_w_lg_w_lg_load_opcode226w227w(i);
	END GENERATE loop21;
	wire_w_lg_w_lg_w_lg_w_lg_do_write58w59w401w402w(0) <= wire_w_lg_w_lg_w_lg_do_write58w59w401w(0) OR wire_w_lg_do_read400w(0);
	wire_w_lg_w_lg_w_lg_rden_wire405w406w407w(0) <= wire_w_lg_w_lg_rden_wire405w406w(0) OR wire_w_lg_stage4_wire404w(0);
	wire_w_lg_w_lg_not_busy397w398w(0) <= wire_w_lg_not_busy397w(0) OR wire_w_lg_addr_overdie395w(0);
	loop22 : FOR i IN 0 TO 22 GENERATE 
		wire_w_lg_w_lg_not_busy389w390w(i) <= wire_w_lg_not_busy389w(i) OR wire_w_lg_stage3_wire387w(i);
	END GENERATE loop22;
	wire_w_lg_w_lg_stage4_wire436w437w(0) <= wire_w_lg_stage4_wire436w(0) OR wire_w_lg_stage3_wire434w(0);
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode229w283w284w285w(0) <= wire_w_lg_w_lg_w_lg_load_opcode229w283w284w(0) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode221w222w223w279w(0);
	loop23 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_load_opcode229w230w231w232w(i) <= wire_w_lg_w_lg_w_lg_load_opcode229w230w231w(i) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode221w222w223w224w(i);
	END GENERATE loop23;
	wire_w_lg_w_lg_w_lg_w_lg_rden_wire405w406w407w408w(0) <= wire_w_lg_w_lg_w_lg_rden_wire405w406w407w(0) OR wire_w_lg_stage3_wire403w(0);
	loop24 : FOR i IN 0 TO 22 GENERATE 
		wire_w_lg_w_lg_w_lg_not_busy389w390w391w(i) <= wire_w_lg_w_lg_not_busy389w390w(i) OR wire_w_lg_addr_overdie385w(i);
	END GENERATE loop24;
	wire_w286w(0) <= wire_w_lg_w_lg_w_lg_w_lg_load_opcode229w283w284w285w(0) OR wire_w_lg_w_lg_load_opcode218w277w(0);
	loop25 : FOR i IN 0 TO 6 GENERATE 
		wire_w233w(i) <= wire_w_lg_w_lg_w_lg_w_lg_load_opcode229w230w231w232w(i) OR wire_w_lg_w_lg_load_opcode218w219w(i);
	END GENERATE loop25;
	wire_w_lg_w286w287w(0) <= wire_w286w(0) OR wire_w_lg_w_lg_load_opcode215w275w(0);
	loop26 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w233w234w(i) <= wire_w233w(i) OR wire_w_lg_w_lg_load_opcode215w216w(i);
	END GENERATE loop26;
	wire_w_lg_w_lg_w286w287w288w(0) <= wire_w_lg_w286w287w(0) OR wire_w273w(0);
	loop27 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w233w234w235w(i) <= wire_w_lg_w233w234w(i) OR wire_w213w(i);
	END GENERATE loop27;
	wire_w_lg_w_lg_w_lg_w286w287w288w289w(0) <= wire_w_lg_w_lg_w286w287w288w(0) OR wire_w271w(0);
	loop28 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w233w234w235w236w(i) <= wire_w_lg_w_lg_w233w234w235w(i) OR wire_w206w(i);
	END GENERATE loop28;
	wire_w_lg_w_lg_w_lg_w_lg_w286w287w288w289w290w(0) <= wire_w_lg_w_lg_w_lg_w286w287w288w289w(0) OR wire_w_lg_w_lg_load_opcode198w269w(0);
	loop29 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_w233w234w235w236w237w(i) <= wire_w_lg_w_lg_w_lg_w233w234w235w236w(i) OR wire_w_lg_w_lg_load_opcode198w199w(i);
	END GENERATE loop29;
	wire_w_lg_w_lg_w_lg_w_lg_w_lg_w286w287w288w289w290w291w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w286w287w288w289w290w(0) OR wire_w_lg_w_lg_load_opcode195w267w(0);
	loop30 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_w_lg_w233w234w235w236w237w238w(i) <= wire_w_lg_w_lg_w_lg_w_lg_w233w234w235w236w237w(i) OR wire_w_lg_w_lg_load_opcode195w196w(i);
	END GENERATE loop30;
	wire_w292w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w_lg_w286w287w288w289w290w291w(0) OR wire_w_lg_w_lg_w_lg_load_opcode185w190w265w(0);
	loop31 : FOR i IN 0 TO 6 GENERATE 
		wire_w239w(i) <= wire_w_lg_w_lg_w_lg_w_lg_w_lg_w233w234w235w236w237w238w(i) OR wire_w_lg_w_lg_w_lg_load_opcode185w190w191w(i);
	END GENERATE loop31;
	wire_w_lg_w292w293w(0) <= wire_w292w(0) OR wire_w_lg_w_lg_w_lg_load_opcode185w186w263w(0);
	loop32 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w239w240w(i) <= wire_w239w(i) OR wire_w_lg_w_lg_w_lg_load_opcode185w186w187w(i);
	END GENERATE loop32;
	wire_w_lg_w_lg_w292w293w294w(0) <= wire_w_lg_w292w293w(0) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode180w181w182w261w(0);
	loop33 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w239w240w241w(i) <= wire_w_lg_w239w240w(i) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode180w181w182w183w(i);
	END GENERATE loop33;
	wire_w_lg_w_lg_w_lg_w292w293w294w295w(0) <= wire_w_lg_w_lg_w292w293w294w(0) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode175w176w177w259w(0);
	loop34 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w239w240w241w242w(i) <= wire_w_lg_w_lg_w239w240w241w(i) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode175w176w177w178w(i);
	END GENERATE loop34;
	wire_w_lg_w_lg_w_lg_w_lg_w292w293w294w295w296w(0) <= wire_w_lg_w_lg_w_lg_w292w293w294w295w(0) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode170w171w172w257w(0);
	loop35 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_w239w240w241w242w243w(i) <= wire_w_lg_w_lg_w_lg_w239w240w241w242w(i) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode170w171w172w173w(i);
	END GENERATE loop35;
	wire_w_lg_w_lg_w_lg_w_lg_w_lg_w292w293w294w295w296w297w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w292w293w294w295w296w(0) OR wire_w_lg_w_lg_load_opcode167w255w(0);
	loop36 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_w_lg_w239w240w241w242w243w244w(i) <= wire_w_lg_w_lg_w_lg_w_lg_w239w240w241w242w243w(i) OR wire_w_lg_w_lg_load_opcode167w168w(i);
	END GENERATE loop36;
	wire_w298w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w_lg_w292w293w294w295w296w297w(0) OR wire_w_lg_w_lg_load_opcode164w253w(0);
	loop37 : FOR i IN 0 TO 6 GENERATE 
		wire_w245w(i) <= wire_w_lg_w_lg_w_lg_w_lg_w_lg_w239w240w241w242w243w244w(i) OR wire_w_lg_w_lg_load_opcode164w165w(i);
	END GENERATE loop37;
	wire_w_lg_w298w299w(0) <= wire_w298w(0) OR wire_w_lg_w_lg_load_opcode159w251w(0);
	loop38 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w245w246w(i) <= wire_w245w(i) OR wire_w_lg_w_lg_load_opcode159w160w(i);
	END GENERATE loop38;
	loop39 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w245w246w247w(i) <= wire_w_lg_w245w246w(i) OR wire_w_lg_shift_opcode155w(i);
	END GENERATE loop39;
	wire_w_lg_w_lg_w137w138w139w(0) <= wire_w_lg_w137w138w(0) OR do_read_nonvolatile;
	wire_w_lg_w137w138w(0) <= wire_w137w(0) OR do_fast_read;
	wire_w_lg_w105w106w(0) <= wire_w105w(0) OR do_ex4baddr;
	wire_w137w(0) <= wire_w_lg_w_lg_w_lg_w_lg_do_read_sid133w134w135w136w(0) OR do_read;
	wire_w105w(0) <= wire_w_lg_w_lg_w_lg_w_lg_do_write58w102w103w104w(0) OR do_4baddr;
	wire_w_lg_w_lg_w_lg_w_lg_do_read400w421w422w423w(0) <= wire_w_lg_w_lg_w_lg_do_read400w421w422w(0) OR do_die_erase;
	wire_w_lg_w_lg_w_lg_w_lg_do_read_sid133w134w135w136w(0) <= wire_w_lg_w_lg_w_lg_do_read_sid133w134w135w(0) OR do_read_rdid;
	wire_w_lg_w_lg_w_lg_w_lg_do_write58w102w103w104w(0) <= wire_w_lg_w_lg_w_lg_do_write58w102w103w(0) OR do_fread_epcq;
	wire_w_lg_w_lg_w_lg_do_read400w421w422w(0) <= wire_w_lg_w_lg_do_read400w421w(0) OR do_sec_erase;
	wire_w_lg_w_lg_w_lg_do_read_sid133w134w135w(0) <= wire_w_lg_w_lg_do_read_sid133w134w(0) OR do_die_erase;
	wire_w_lg_w_lg_w_lg_do_read_stat431w432w433w(0) <= wire_w_lg_w_lg_do_read_stat431w432w(0) OR do_read_nonvolatile;
	wire_w_lg_w_lg_w_lg_do_write58w102w103w(0) <= wire_w_lg_w_lg_do_write58w102w(0) OR do_die_erase;
	wire_w_lg_w_lg_do_read400w435w(0) <= wire_w_lg_do_read400w(0) OR do_read_sid;
	wire_w_lg_w_lg_do_read400w421w(0) <= wire_w_lg_do_read400w(0) OR do_write;
	wire_w_lg_w_lg_do_read_sid133w134w(0) <= wire_w_lg_do_read_sid133w(0) OR do_sec_erase;
	wire_w_lg_w_lg_do_read_stat431w432w(0) <= wire_w_lg_do_read_stat431w(0) OR do_read_volatile;
	wire_w_lg_w_lg_do_write58w102w(0) <= wire_w_lg_do_write58w(0) OR do_bulk_erase;
	wire_w_lg_w_lg_do_write58w59w(0) <= wire_w_lg_do_write58w(0) OR do_die_erase;
	wire_w_lg_data0out_wire439w(0) <= data0out_wire OR wire_w_dataout_wire_range438w(0);
	wire_w_lg_do_4baddr334w(0) <= do_4baddr OR wire_w_lg_do_ex4baddr333w(0);
	wire_w_lg_do_ex4baddr333w(0) <= do_ex4baddr OR wire_w_lg_do_bulk_erase332w(0);
	wire_w_lg_do_read400w(0) <= do_read OR do_fast_read;
	wire_w_lg_do_read_rdid111w(0) <= do_read_rdid OR wire_w_lg_w_lg_do_read_stat109w110w(0);
	wire_w_lg_do_read_sid133w(0) <= do_read_sid OR do_write;
	wire_w_lg_do_read_stat431w(0) <= do_read_stat OR do_read_rdid;
	wire_w_lg_do_sec_erase40w(0) <= do_sec_erase OR do_die_erase;
	wire_w_lg_do_wren335w(0) <= do_wren OR wire_w_lg_do_4baddr334w(0);
	wire_w_lg_do_write58w(0) <= do_write OR do_sec_erase;
	wire_w_lg_load_opcode301w(0) <= load_opcode OR shift_opcode;
	wire_w_lg_rden_wire405w(0) <= rden_wire OR wren_wire;
	add_rollover <= add_rollover_reg;
	addr_overdie <= '0';
	addr_overdie_pos <= '0';
	addr_reg_overdie <= (OTHERS => '0');
	b4addr_opcode <= (OTHERS => '0');
	berase_opcode <= (OTHERS => '0');
	busy <= busy_wire;
	busy_wire <= ((((((((((((((do_read_rdid OR do_read_sid) OR do_read) OR do_fast_read) OR do_write) OR do_sec_prot) OR do_read_stat) OR do_sec_erase) OR do_bulk_erase) OR do_die_erase) OR do_4baddr) OR do_read_volatile) OR do_fread_epcq) OR do_read_nonvolatile) OR do_ex4baddr);
	clkin_wire <= clkin;
	clr_addmsb_wire <= ((wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range89w94w413w414w(0) OR wire_w_lg_w_lg_w_lg_do_read352w353w412w(0)) OR wire_w_lg_w_lg_w_lg_w_lg_do_sec_erase40w409w410w411w(0));
	clr_endrbyte_wire <= ((((wire_w_lg_do_read400w(0) AND (NOT wire_gen_cntr_q(2))) AND wire_gen_cntr_q(1)) AND wire_gen_cntr_q(0)) OR clr_read_wire2);
	clr_read_wire <= clr_read_reg;
	clr_read_wire2 <= clr_read_reg2;
	clr_write_wire2 <= '0';
	data0out_wire <= wire_arriav_asmiblock2_data1in;
	data_valid <= data_valid_wire;
	data_valid_wire <= dvalid_reg2;
	dataoe_wire <= ( "1" & "1" & "0" & "1");
	dataout <= ( read_data_reg(7 DOWNTO 0));
	dataout_wire <= ( "0000");
	derase_opcode <= (OTHERS => '0');
	do_4baddr <= '0';
	do_bulk_erase <= '0';
	do_die_erase <= '0';
	do_ex4baddr <= '0';
	do_fast_read <= '0';
	do_fread_epcq <= '0';
	do_freadwrv_polling <= '0';
	do_memadd <= '0';
	do_polling <= ((do_write_polling OR do_sprot_polling) OR do_freadwrv_polling);
	do_read <= (((wire_w_lg_read_rdid_wire7w(0) AND wire_w_lg_read_sid_wire6w(0)) AND wire_w_lg_sec_protect_wire5w(0)) AND read_wire);
	do_read_nonvolatile <= '0';
	do_read_rdid <= '0';
	do_read_sid <= '0';
	do_read_stat <= '0';
	do_read_volatile <= '0';
	do_sec_erase <= '0';
	do_sec_prot <= '0';
	do_sprot_polling <= '0';
	do_wait_dummyclk <= '0';
	do_wren <= '0';
	do_write <= '0';
	do_write_polling <= '0';
	do_write_volatile <= '0';
	end1_cyc_gen_cntr_wire <= (wire_gen_cntr_w_lg_w_q_range99w100w(0) AND (NOT wire_gen_cntr_q(0)));
	end1_cyc_normal_in_wire <= ((((((((((wire_stage_cntr_w_lg_w_lg_w_q_range88w93w119w(0) AND (NOT wire_gen_cntr_q(2))) AND wire_gen_cntr_q(1)) AND wire_gen_cntr_q(0)) OR wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range88w93w119w120w121w(0)) OR (do_read AND end_read)) OR (do_fast_read AND end_fast_read)) OR wire_w_lg_w_lg_w_lg_w_lg_do_write58w102w103w116w(0)) OR wire_w_lg_do_write56w(0)) OR ((do_read_stat AND start_poll) AND wire_w_lg_st_busy_wire113w(0))) OR wire_w_lg_w_lg_do_read_rdid111w112w(0));
	end1_cyc_reg_in_wire <= end1_cyc_normal_in_wire;
	end_add_cycle <= wire_mux211_dataout;
	end_add_cycle_mux_datab_wire <= (wire_addbyte_cntr_q(2) AND wire_addbyte_cntr_q(1));
	end_fast_read <= end_read_reg;
	end_one_cyc_pos <= end1_cyc_reg2;
	end_one_cycle <= end1_cyc_reg;
	end_op_wire <= (((((((((((wire_stage_cntr_w_lg_w_q_range89w94w(0) AND ((wire_w_lg_w_lg_w_lg_w_lg_do_read352w353w354w355w(0) OR (do_read AND end_read)) OR (do_fast_read AND end_fast_read))) OR (wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range89w92w347w348w(0) AND wire_w_lg_do_polling189w(0))) OR ((((((do_read_rdid AND end_one_cyc_pos) AND wire_stage_cntr_q(1)) AND wire_stage_cntr_q(0)) AND wire_addbyte_cntr_q(2)) AND wire_addbyte_cntr_q(1)) AND wire_addbyte_cntr_w_lg_w_q_range147w148w(0))) OR (wire_w_lg_w_lg_start_poll338w339w(0) AND wire_w_lg_st_busy_wire113w(0))) OR wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range89w90w91w336w337w(0)) OR wire_w_lg_w_lg_w_lg_w_lg_do_write58w102w103w116w(0)) OR wire_w_lg_w_lg_do_write49w331w(0)) OR wire_w_lg_do_write56w(0)) OR wire_stage_cntr_w330w(0)) OR wire_stage_cntr_w_lg_w325w326w(0)) OR (wire_stage_cntr_w_lg_w_lg_w_q_range89w92w320w(0) AND ((do_write_volatile OR do_read_volatile) OR wire_w_lg_do_read_nonvolatile318w(0))));
	end_operation <= end_op_reg;
	end_ophdly <= end_op_hdlyreg;
	end_pgwr_data <= '0';
	end_read <= end_read_reg;
	end_read_byte <= (end_rbyte_reg AND wire_w_lg_addr_overdie499w(0));
	exb4addr_opcode <= (OTHERS => '0');
	fast_read_opcode <= (OTHERS => '0');
	freadwrv_sdoin <= '0';
	in_operation <= busy_wire;
	load_opcode <= ((((wire_stage_cntr_w_lg_w_q_range89w90w(0) AND wire_stage_cntr_w_lg_w_q_range88w93w(0)) AND (NOT wire_gen_cntr_q(2))) AND wire_gen_cntr_w_lg_w_q_range97w98w(0)) AND wire_gen_cntr_q(0));
	memadd_sdoin <= add_msb_reg;
	ncs_reg_ena_wire <= (((wire_stage_cntr_w_lg_w_lg_w_q_range89w90w91w(0) AND end_one_cyc_pos) OR addr_overdie_pos) OR end_operation);
	not_busy <= busy_det_reg;
	oe_wire <= '0';
	pagewr_buf_not_empty <= ( "1");
	rden_wire <= rden;
	rdid_opcode <= (OTHERS => '0');
	rdummyclk_opcode <= (OTHERS => '0');
	read_address <= ( read_add_reg(23 DOWNTO 0));
	read_data_reg_in_wire <= ( read_dout_reg(7 DOWNTO 0));
	read_opcode <= "00000011";
	read_rdid_wire <= '0';
	read_sid_wire <= '0';
	read_wire <= read_reg;
	rflagstat_opcode <= (OTHERS => '0');
	rnvdummyclk_opcode <= (OTHERS => '0');
	rsid_opcode <= (OTHERS => '0');
	rsid_sdoin <= '0';
	rstat_opcode <= (OTHERS => '0');
	scein_wire <= wire_ncs_reg_w_lg_q373w(0);
	sdoin_wire <= to_sdoin_wire;
	sec_protect_wire <= '0';
	secprot_opcode <= (OTHERS => '0');
	secprot_sdoin <= '0';
	serase_opcode <= (OTHERS => '0');
	shift_opcode <= shift_op_reg;
	shift_opdata <= stage2_wire;
	shift_pgwr_data <= '0';
	st_busy_wire <= '0';
	stage2_wire <= stage2_reg;
	stage3_wire <= stage3_reg;
	stage4_wire <= stage4_reg;
	start_frpoll <= '0';
	start_poll <= ((start_wrpoll OR start_sppoll) OR start_frpoll);
	start_sppoll <= '0';
	start_wrpoll <= '0';
	to_sdoin_wire <= ((((((shift_opdata AND asmi_opcode_reg(7)) OR rsid_sdoin) OR memadd_sdoin) OR write_sdoin) OR secprot_sdoin) OR freadwrv_sdoin);
	wren_opcode <= (OTHERS => '0');
	wren_wire <= '1';
	write_opcode <= (OTHERS => '0');
	write_prot_true <= '0';
	write_sdoin <= '0';
	wrvolatile_opcode <= (OTHERS => '0');
	wire_w_addr_range396w(0) <= addr(0);
	wire_w_addr_range388w <= addr(23 DOWNTO 1);
	wire_w_addr_reg_overdie_range394w(0) <= addr_reg_overdie(0);
	wire_w_addr_reg_overdie_range384w <= addr_reg_overdie(23 DOWNTO 1);
	wire_w_b4addr_opcode_range252w(0) <= b4addr_opcode(0);
	wire_w_b4addr_opcode_range161w <= b4addr_opcode(7 DOWNTO 1);
	wire_w_berase_opcode_range256w(0) <= berase_opcode(0);
	wire_w_berase_opcode_range169w <= berase_opcode(7 DOWNTO 1);
	wire_w_dataout_wire_range438w(0) <= dataout_wire(1);
	wire_w_derase_opcode_range258w(0) <= derase_opcode(0);
	wire_w_derase_opcode_range174w <= derase_opcode(7 DOWNTO 1);
	wire_w_exb4addr_opcode_range250w(0) <= exb4addr_opcode(0);
	wire_w_exb4addr_opcode_range156w <= exb4addr_opcode(7 DOWNTO 1);
	wire_w_fast_read_opcode_range274w(0) <= fast_read_opcode(0);
	wire_w_fast_read_opcode_range214w <= fast_read_opcode(7 DOWNTO 1);
	wire_w_pagewr_buf_not_empty_range54w(0) <= pagewr_buf_not_empty(0);
	wire_w_rdid_opcode_range280w(0) <= rdid_opcode(0);
	wire_w_rdid_opcode_range225w <= rdid_opcode(7 DOWNTO 1);
	wire_w_rdummyclk_opcode_range272w(0) <= rdummyclk_opcode(0);
	wire_w_rdummyclk_opcode_range207w <= rdummyclk_opcode(7 DOWNTO 1);
	wire_w_read_opcode_range276w(0) <= read_opcode(0);
	wire_w_read_opcode_range217w <= read_opcode(7 DOWNTO 1);
	wire_w_rflagstat_opcode_range262w(0) <= rflagstat_opcode(0);
	wire_w_rflagstat_opcode_range184w <= rflagstat_opcode(7 DOWNTO 1);
	wire_w_rnvdummyclk_opcode_range268w(0) <= rnvdummyclk_opcode(0);
	wire_w_rnvdummyclk_opcode_range197w <= rnvdummyclk_opcode(7 DOWNTO 1);
	wire_w_rsid_opcode_range282w(0) <= rsid_opcode(0);
	wire_w_rsid_opcode_range228w <= rsid_opcode(7 DOWNTO 1);
	wire_w_rstat_opcode_range264w(0) <= rstat_opcode(0);
	wire_w_rstat_opcode_range188w <= rstat_opcode(7 DOWNTO 1);
	wire_w_secprot_opcode_range278w(0) <= secprot_opcode(0);
	wire_w_secprot_opcode_range220w <= secprot_opcode(7 DOWNTO 1);
	wire_w_serase_opcode_range260w(0) <= serase_opcode(0);
	wire_w_serase_opcode_range179w <= serase_opcode(7 DOWNTO 1);
	wire_w_wren_opcode_range254w(0) <= wren_opcode(0);
	wire_w_wren_opcode_range166w <= wren_opcode(7 DOWNTO 1);
	wire_w_write_opcode_range266w(0) <= write_opcode(0);
	wire_w_write_opcode_range192w <= write_opcode(7 DOWNTO 1);
	wire_w_wrvolatile_opcode_range270w(0) <= wrvolatile_opcode(0);
	wire_w_wrvolatile_opcode_range200w <= wrvolatile_opcode(7 DOWNTO 1);
	wire_addbyte_cntr_w_lg_w_q_range144w149w(0) <= wire_addbyte_cntr_w_q_range144w(0) AND wire_addbyte_cntr_w_lg_w_q_range147w148w(0);
	wire_addbyte_cntr_w_lg_w_q_range147w148w(0) <= NOT wire_addbyte_cntr_w_q_range147w(0);
	wire_addbyte_cntr_clk_en <= wire_stage_cntr_w143w(0);
	wire_stage_cntr_w143w(0) <= ((wire_stage_cntr_w_lg_w_lg_w_q_range89w92w140w(0) AND wire_w_lg_w_lg_w137w138w139w(0)) OR addr_overdie) OR end_operation;
	wire_addbyte_cntr_clock <= wire_w_lg_clkin_wire87w(0);
	wire_addbyte_cntr_sclr <= wire_w_lg_end_operation86w(0);
	wire_w_lg_end_operation86w(0) <= end_operation OR addr_overdie;
	wire_addbyte_cntr_w_q_range147w(0) <= wire_addbyte_cntr_q(0);
	wire_addbyte_cntr_w_q_range144w(0) <= wire_addbyte_cntr_q(1);
	addbyte_cntr :  a_graycounter
	  GENERIC MAP (
		WIDTH => 3
	  )
	  PORT MAP ( 
		aclr => reset,
		clk_en => wire_addbyte_cntr_clk_en,
		clock => wire_addbyte_cntr_clock,
		q => wire_addbyte_cntr_q,
		sclr => wire_addbyte_cntr_sclr
	  );
	wire_gen_cntr_w_lg_w_q_range99w100w(0) <= wire_gen_cntr_w_q_range99w(0) AND wire_gen_cntr_w_lg_w_q_range97w98w(0);
	wire_gen_cntr_w_lg_w_q_range97w98w(0) <= NOT wire_gen_cntr_w_q_range97w(0);
	wire_gen_cntr_clk_en <= wire_w_lg_w_lg_w_lg_in_operation26w27w28w(0);
	wire_w_lg_w_lg_w_lg_in_operation26w27w28w(0) <= ((in_operation AND wire_w_lg_end_ophdly25w(0)) OR do_wait_dummyclk) OR addr_overdie;
	wire_gen_cntr_sclr <= wire_w_lg_w_lg_end1_cyc_reg_in_wire29w30w(0);
	wire_w_lg_w_lg_end1_cyc_reg_in_wire29w30w(0) <= (end1_cyc_reg_in_wire OR addr_overdie) OR do_wait_dummyclk;
	wire_gen_cntr_w_q_range97w(0) <= wire_gen_cntr_q(1);
	wire_gen_cntr_w_q_range99w(0) <= wire_gen_cntr_q(2);
	gen_cntr :  a_graycounter
	  GENERIC MAP (
		WIDTH => 3
	  )
	  PORT MAP ( 
		aclr => reset,
		clk_en => wire_gen_cntr_clk_en,
		clock => clkin_wire,
		q => wire_gen_cntr_q,
		sclr => wire_gen_cntr_sclr
	  );
	wire_stage_cntr_w_lg_w325w326w(0) <= wire_stage_cntr_w325w(0) AND end_one_cycle;
	wire_stage_cntr_w325w(0) <= wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range89w92w322w323w324w(0) AND end_add_cycle;
	wire_stage_cntr_w330w(0) <= wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range89w92w327w328w329w(0) AND end_one_cycle;
	wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range89w92w322w323w324w(0) <= wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range89w92w322w323w(0) AND wire_w_lg_do_read_stat38w(0);
	wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range89w92w327w328w329w(0) <= wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range89w92w327w328w(0) AND wire_w_lg_do_read_stat38w(0);
	wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range89w90w91w336w337w(0) <= wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range89w90w91w336w(0) AND end_one_cycle;
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range89w94w413w414w(0) <= wire_stage_cntr_w_lg_w_lg_w_q_range89w94w413w(0) AND end_one_cyc_pos;
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range89w92w322w323w(0) <= wire_stage_cntr_w_lg_w_lg_w_q_range89w92w322w(0) AND wire_w_lg_do_wren39w(0);
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range89w92w347w348w(0) <= wire_stage_cntr_w_lg_w_lg_w_q_range89w92w347w(0) AND end_one_cycle;
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range89w92w327w328w(0) <= wire_stage_cntr_w_lg_w_lg_w_q_range89w92w327w(0) AND wire_w_lg_do_wren39w(0);
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range89w90w91w336w(0) <= wire_stage_cntr_w_lg_w_lg_w_q_range89w90w91w(0) AND wire_w_lg_do_wren335w(0);
	wire_stage_cntr_w_lg_w_lg_w_q_range89w94w413w(0) <= wire_stage_cntr_w_lg_w_q_range89w94w(0) AND end_add_cycle;
	wire_stage_cntr_w_lg_w_lg_w_q_range89w92w322w(0) <= wire_stage_cntr_w_lg_w_q_range89w92w(0) AND wire_w_lg_do_sec_erase40w(0);
	wire_stage_cntr_w_lg_w_lg_w_q_range89w92w347w(0) <= wire_stage_cntr_w_lg_w_q_range89w92w(0) AND do_read_stat;
	wire_stage_cntr_w_lg_w_lg_w_q_range89w92w327w(0) <= wire_stage_cntr_w_lg_w_q_range89w92w(0) AND do_sec_prot;
	wire_stage_cntr_w_lg_w_lg_w_q_range89w92w140w(0) <= wire_stage_cntr_w_lg_w_q_range89w92w(0) AND end_one_cyc_pos;
	wire_stage_cntr_w_lg_w_lg_w_q_range89w92w320w(0) <= wire_stage_cntr_w_lg_w_q_range89w92w(0) AND end_one_cycle;
	wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range88w93w119w120w121w(0) <= wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range88w93w119w120w(0) AND end1_cyc_gen_cntr_wire;
	wire_stage_cntr_w_lg_w_lg_w_q_range88w93w119w(0) <= wire_stage_cntr_w_lg_w_q_range88w93w(0) AND wire_stage_cntr_w_lg_w_q_range89w90w(0);
	wire_stage_cntr_w_lg_w_lg_w_q_range89w90w91w(0) <= wire_stage_cntr_w_lg_w_q_range89w90w(0) AND wire_stage_cntr_w_q_range88w(0);
	wire_stage_cntr_w_lg_w_q_range89w94w(0) <= wire_stage_cntr_w_q_range89w(0) AND wire_stage_cntr_w_lg_w_q_range88w93w(0);
	wire_stage_cntr_w_lg_w_q_range89w92w(0) <= wire_stage_cntr_w_q_range89w(0) AND wire_stage_cntr_w_q_range88w(0);
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range88w93w119w120w(0) <= NOT wire_stage_cntr_w_lg_w_lg_w_q_range88w93w119w(0);
	wire_stage_cntr_w_lg_w_q_range88w93w(0) <= NOT wire_stage_cntr_w_q_range88w(0);
	wire_stage_cntr_w_lg_w_q_range89w90w(0) <= NOT wire_stage_cntr_w_q_range89w(0);
	wire_stage_cntr_clk_en <= wire_w_lg_w_lg_w_lg_w82w83w84w85w(0);
	wire_w_lg_w_lg_w_lg_w82w83w84w85w(0) <= (((((((((((((in_operation AND end_one_cycle) AND (NOT (stage3_wire AND wire_w_lg_end_add_cycle69w(0)))) AND (NOT (stage4_wire AND wire_w_lg_end_read66w(0)))) AND (NOT (stage4_wire AND wire_w_lg_end_fast_read63w(0)))) AND (NOT ((wire_w_lg_w_lg_do_write58w59w(0) OR do_bulk_erase) AND write_prot_true))) AND (NOT wire_w_lg_do_write56w(0))) AND (NOT (stage3_wire AND st_busy_wire))) AND (NOT (wire_w_lg_do_write49w(0) AND wire_w_lg_end_pgwr_data48w(0)))) AND (NOT (stage2_wire AND do_wren))) AND (NOT (((wire_w_lg_stage3_wire41w(0) AND wire_w_lg_do_wren39w(0)) AND wire_w_lg_do_read_stat38w(0)) AND wire_w_lg_do_read_rdid37w(0)))) AND (NOT (stage3_wire AND ((do_write_volatile OR do_read_volatile) OR do_read_nonvolatile)))) OR wire_w_lg_w_lg_stage3_wire31w32w(0)) OR addr_overdie) OR end_ophdly;
	wire_stage_cntr_sclr <= wire_w_lg_end_operation86w(0);
	wire_stage_cntr_w_q_range88w(0) <= wire_stage_cntr_q(0);
	wire_stage_cntr_w_q_range89w(0) <= wire_stage_cntr_q(1);
	stage_cntr :  a_graycounter
	  GENERIC MAP (
		WIDTH => 2
	  )
	  PORT MAP ( 
		aclr => reset,
		clk_en => wire_stage_cntr_clk_en,
		clock => clkin_wire,
		q => wire_stage_cntr_q,
		sclr => wire_stage_cntr_sclr
	  );
	arriav_asmiblock2 :  cyclonev_asmiblock
	  PORT MAP ( 
		data0oe => dataoe_wire(0),
		data0out => sdoin_wire,
		data1in => wire_arriav_asmiblock2_data1in,
		data1oe => dataoe_wire(1),
		data2oe => dataoe_wire(2),
		data2out => wire_vcc,
		data3oe => dataoe_wire(3),
		data3out => wire_vcc,
		dclk => clkin_wire,
		oe => oe_wire,
		sce => scein_wire
	  );
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN add_msb_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_add_msb_reg_ena = '1') THEN 
				IF (clr_addmsb_wire = '1') THEN add_msb_reg <= '0';
				ELSE add_msb_reg <= addr_reg(23);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_add_msb_reg_ena <= ((((wire_w_lg_w_lg_w_lg_w_lg_do_read400w421w422w423w(0) AND (NOT (wire_w_lg_w_lg_do_write58w59w(0) AND wire_w_lg_do_memadd418w(0)))) AND wire_stage_cntr_q(1)) AND wire_stage_cntr_q(0)) OR clr_addmsb_wire);
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN add_rollover_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN add_rollover_reg <= (wire_read_add_cntr_q(23) OR clr_read_wire2);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(0) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(0) = '1') THEN addr_reg(0) <= wire_addr_reg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(1) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(1) = '1') THEN addr_reg(1) <= wire_addr_reg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(2) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(2) = '1') THEN addr_reg(2) <= wire_addr_reg_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(3) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(3) = '1') THEN addr_reg(3) <= wire_addr_reg_d(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(4) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(4) = '1') THEN addr_reg(4) <= wire_addr_reg_d(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(5) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(5) = '1') THEN addr_reg(5) <= wire_addr_reg_d(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(6) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(6) = '1') THEN addr_reg(6) <= wire_addr_reg_d(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(7) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(7) = '1') THEN addr_reg(7) <= wire_addr_reg_d(7);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(8) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(8) = '1') THEN addr_reg(8) <= wire_addr_reg_d(8);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(9) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(9) = '1') THEN addr_reg(9) <= wire_addr_reg_d(9);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(10) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(10) = '1') THEN addr_reg(10) <= wire_addr_reg_d(10);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(11) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(11) = '1') THEN addr_reg(11) <= wire_addr_reg_d(11);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(12) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(12) = '1') THEN addr_reg(12) <= wire_addr_reg_d(12);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(13) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(13) = '1') THEN addr_reg(13) <= wire_addr_reg_d(13);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(14) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(14) = '1') THEN addr_reg(14) <= wire_addr_reg_d(14);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(15) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(15) = '1') THEN addr_reg(15) <= wire_addr_reg_d(15);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(16) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(16) = '1') THEN addr_reg(16) <= wire_addr_reg_d(16);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(17) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(17) = '1') THEN addr_reg(17) <= wire_addr_reg_d(17);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(18) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(18) = '1') THEN addr_reg(18) <= wire_addr_reg_d(18);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(19) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(19) = '1') THEN addr_reg(19) <= wire_addr_reg_d(19);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(20) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(20) = '1') THEN addr_reg(20) <= wire_addr_reg_d(20);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(21) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(21) = '1') THEN addr_reg(21) <= wire_addr_reg_d(21);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(22) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(22) = '1') THEN addr_reg(22) <= wire_addr_reg_d(22);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(23) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(23) = '1') THEN addr_reg(23) <= wire_addr_reg_d(23);
			END IF;
		END IF;
	END PROCESS;
	wire_addr_reg_d <= ( wire_w_lg_w_lg_w_lg_not_busy389w390w391w & wire_w_lg_w_lg_not_busy397w398w);
	loop40 : FOR i IN 0 TO 23 GENERATE
		wire_addr_reg_ena(i) <= wire_w_lg_w_lg_w_lg_w_lg_rden_wire405w406w407w408w(0);
	END GENERATE loop40;
	wire_addr_reg_w_q_range386w <= addr_reg(22 DOWNTO 0);
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN asmi_opcode_reg(0) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(0) = '1') THEN asmi_opcode_reg(0) <= wire_asmi_opcode_reg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN asmi_opcode_reg(1) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(1) = '1') THEN asmi_opcode_reg(1) <= wire_asmi_opcode_reg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN asmi_opcode_reg(2) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(2) = '1') THEN asmi_opcode_reg(2) <= wire_asmi_opcode_reg_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN asmi_opcode_reg(3) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(3) = '1') THEN asmi_opcode_reg(3) <= wire_asmi_opcode_reg_d(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN asmi_opcode_reg(4) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(4) = '1') THEN asmi_opcode_reg(4) <= wire_asmi_opcode_reg_d(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN asmi_opcode_reg(5) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(5) = '1') THEN asmi_opcode_reg(5) <= wire_asmi_opcode_reg_d(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN asmi_opcode_reg(6) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(6) = '1') THEN asmi_opcode_reg(6) <= wire_asmi_opcode_reg_d(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN asmi_opcode_reg(7) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(7) = '1') THEN asmi_opcode_reg(7) <= wire_asmi_opcode_reg_d(7);
			END IF;
		END IF;
	END PROCESS;
	wire_asmi_opcode_reg_d <= ( wire_w_lg_w_lg_w245w246w247w & wire_w_lg_w298w299w);
	loop41 : FOR i IN 0 TO 7 GENERATE
		wire_asmi_opcode_reg_ena(i) <= wire_w_lg_load_opcode301w(0);
	END GENERATE loop41;
	wire_asmi_opcode_reg_w_q_range154w <= asmi_opcode_reg(6 DOWNTO 0);
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN busy_det_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN busy_det_reg <= wire_w_lg_busy_wire1w(0);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN clr_read_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN clr_read_reg <= ((do_read_sid OR do_sec_prot) OR end_operation);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN clr_read_reg2 <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN clr_read_reg2 <= clr_read_reg;
		END IF;
	END PROCESS;
	dffe3 <= '0';
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN dvalid_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_dvalid_reg_ena = '1') THEN 
				IF (wire_dvalid_reg_sclr = '1') THEN dvalid_reg <= '0';
				ELSE dvalid_reg <= wire_w_lg_end_read_byte474w(0);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_dvalid_reg_ena <= wire_w_lg_do_read400w(0);
	wire_dvalid_reg_sclr <= (end_op_wire OR end_operation);
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN dvalid_reg2 <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN dvalid_reg2 <= dvalid_reg;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN end1_cyc_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN end1_cyc_reg <= end1_cyc_reg_in_wire;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN end1_cyc_reg2 <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN end1_cyc_reg2 <= end_one_cycle;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN end_op_hdlyreg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN end_op_hdlyreg <= end_operation;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN end_op_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN end_op_reg <= end_op_wire;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN end_rbyte_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_end_rbyte_reg_ena = '1') THEN 
				IF (wire_end_rbyte_reg_sclr = '1') THEN end_rbyte_reg <= '0';
				ELSE end_rbyte_reg <= wire_w_lg_w_lg_w_lg_do_read400w467w468w(0);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_end_rbyte_reg_ena <= ((wire_gen_cntr_w_lg_w_q_range99w100w(0) AND wire_gen_cntr_q(0)) OR clr_endrbyte_wire);
	wire_end_rbyte_reg_sclr <= (clr_endrbyte_wire OR addr_overdie);
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN end_read_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN end_read_reg <= (((wire_w_lg_rden_wire501w(0) AND wire_w_lg_do_read400w(0)) AND data_valid_wire) AND end_read_byte);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN ncs_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (ncs_reg_ena_wire = '1') THEN 
				IF (wire_ncs_reg_sclr = '1') THEN ncs_reg <= '0';
				ELSE ncs_reg <= '1';
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_ncs_reg_sclr <= (end_operation OR addr_overdie_pos);
	wire_ncs_reg_w_lg_q373w(0) <= NOT ncs_reg;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(0) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(0) = '1') THEN read_add_reg(0) <= wire_read_add_reg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(1) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(1) = '1') THEN read_add_reg(1) <= wire_read_add_reg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(2) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(2) = '1') THEN read_add_reg(2) <= wire_read_add_reg_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(3) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(3) = '1') THEN read_add_reg(3) <= wire_read_add_reg_d(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(4) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(4) = '1') THEN read_add_reg(4) <= wire_read_add_reg_d(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(5) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(5) = '1') THEN read_add_reg(5) <= wire_read_add_reg_d(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(6) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(6) = '1') THEN read_add_reg(6) <= wire_read_add_reg_d(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(7) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(7) = '1') THEN read_add_reg(7) <= wire_read_add_reg_d(7);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(8) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(8) = '1') THEN read_add_reg(8) <= wire_read_add_reg_d(8);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(9) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(9) = '1') THEN read_add_reg(9) <= wire_read_add_reg_d(9);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(10) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(10) = '1') THEN read_add_reg(10) <= wire_read_add_reg_d(10);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(11) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(11) = '1') THEN read_add_reg(11) <= wire_read_add_reg_d(11);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(12) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(12) = '1') THEN read_add_reg(12) <= wire_read_add_reg_d(12);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(13) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(13) = '1') THEN read_add_reg(13) <= wire_read_add_reg_d(13);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(14) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(14) = '1') THEN read_add_reg(14) <= wire_read_add_reg_d(14);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(15) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(15) = '1') THEN read_add_reg(15) <= wire_read_add_reg_d(15);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(16) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(16) = '1') THEN read_add_reg(16) <= wire_read_add_reg_d(16);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(17) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(17) = '1') THEN read_add_reg(17) <= wire_read_add_reg_d(17);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(18) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(18) = '1') THEN read_add_reg(18) <= wire_read_add_reg_d(18);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(19) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(19) = '1') THEN read_add_reg(19) <= wire_read_add_reg_d(19);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(20) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(20) = '1') THEN read_add_reg(20) <= wire_read_add_reg_d(20);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(21) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(21) = '1') THEN read_add_reg(21) <= wire_read_add_reg_d(21);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(22) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(22) = '1') THEN read_add_reg(22) <= wire_read_add_reg_d(22);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_add_reg(23) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_add_reg_ena(23) = '1') THEN read_add_reg(23) <= wire_read_add_reg_d(23);
			END IF;
		END IF;
	END PROCESS;
	wire_read_add_reg_d <= ( wire_read_add_cntr_q(23 DOWNTO 0));
	loop42 : FOR i IN 0 TO 23 GENERATE
		wire_read_add_reg_ena(i) <= wire_w_lg_w_lg_end_read_byte474w486w(0);
	END GENERATE loop42;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_data_reg(0) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(0) = '1') THEN read_data_reg(0) <= wire_read_data_reg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_data_reg(1) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(1) = '1') THEN read_data_reg(1) <= wire_read_data_reg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_data_reg(2) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(2) = '1') THEN read_data_reg(2) <= wire_read_data_reg_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_data_reg(3) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(3) = '1') THEN read_data_reg(3) <= wire_read_data_reg_d(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_data_reg(4) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(4) = '1') THEN read_data_reg(4) <= wire_read_data_reg_d(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_data_reg(5) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(5) = '1') THEN read_data_reg(5) <= wire_read_data_reg_d(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_data_reg(6) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(6) = '1') THEN read_data_reg(6) <= wire_read_data_reg_d(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_data_reg(7) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(7) = '1') THEN read_data_reg(7) <= wire_read_data_reg_d(7);
			END IF;
		END IF;
	END PROCESS;
	wire_read_data_reg_d <= ( read_data_reg_in_wire(7 DOWNTO 0));
	loop43 : FOR i IN 0 TO 7 GENERATE
		wire_read_data_reg_ena(i) <= wire_w470w(0);
	END GENERATE loop43;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_dout_reg(0) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(0) = '1') THEN read_dout_reg(0) <= wire_read_dout_reg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_dout_reg(1) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(1) = '1') THEN read_dout_reg(1) <= wire_read_dout_reg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_dout_reg(2) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(2) = '1') THEN read_dout_reg(2) <= wire_read_dout_reg_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_dout_reg(3) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(3) = '1') THEN read_dout_reg(3) <= wire_read_dout_reg_d(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_dout_reg(4) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(4) = '1') THEN read_dout_reg(4) <= wire_read_dout_reg_d(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_dout_reg(5) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(5) = '1') THEN read_dout_reg(5) <= wire_read_dout_reg_d(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_dout_reg(6) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(6) = '1') THEN read_dout_reg(6) <= wire_read_dout_reg_d(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_dout_reg(7) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(7) = '1') THEN read_dout_reg(7) <= wire_read_dout_reg_d(7);
			END IF;
		END IF;
	END PROCESS;
	wire_read_dout_reg_d <= ( read_dout_reg(6 DOWNTO 0) & wire_w_lg_data0out_wire439w);
	loop44 : FOR i IN 0 TO 7 GENERATE
		wire_read_dout_reg_ena(i) <= wire_w_lg_w_lg_stage4_wire436w437w(0);
	END GENERATE loop44;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_reg_ena = '1') THEN 
				IF (clr_read_wire = '1') THEN read_reg <= '0';
				ELSE read_reg <= read;
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_read_reg_ena <= ((wire_w_lg_busy_wire1w(0) AND rden_wire) OR clr_read_wire);
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN shift_op_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN shift_op_reg <= wire_stage_cntr_w_lg_w_lg_w_q_range89w90w91w(0);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN stage2_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN stage2_reg <= wire_stage_cntr_w_lg_w_lg_w_q_range89w90w91w(0);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN stage3_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN stage3_reg <= wire_stage_cntr_w_lg_w_q_range89w92w(0);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN stage4_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN stage4_reg <= wire_stage_cntr_w_lg_w_q_range89w94w(0);
		END IF;
	END PROCESS;
	wire_read_add_cntr_clk_en <= wire_w_lg_w_lg_w_lg_rden_wire476w477w478w(0);
	wire_w_lg_w_lg_w_lg_rden_wire476w477w478w(0) <= ((rden_wire AND not_busy) OR data_valid_wire) OR add_rollover;
	wire_read_add_cntr_data <= ( "0" & addr(23 DOWNTO 0));
	wire_read_add_cntr_sload <= wire_w_lg_rden_wire476w(0);
	wire_w_lg_rden_wire476w(0) <= rden_wire AND not_busy;
	read_add_cntr :  lpm_counter
	  GENERIC MAP (
		lpm_direction => "UP",
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 25
	  )
	  PORT MAP ( 
		aclr => reset,
		clk_en => wire_read_add_cntr_clk_en,
		clock => clkin_wire,
		data => wire_read_add_cntr_data,
		q => wire_read_add_cntr_q,
		sclr => add_rollover,
		sload => wire_read_add_cntr_sload
	  );
	wire_mux211_dataout <= end_add_cycle_mux_datab_wire WHEN do_fast_read = '1'  ELSE wire_addbyte_cntr_w_lg_w_q_range144w149w(0);

 END RTL; --asmicont_altasmi_parallel_qth2
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY asmicont IS
	PORT
	(
		addr		: IN STD_LOGIC_VECTOR (23 DOWNTO 0);
		clkin		: IN STD_LOGIC ;
		rden		: IN STD_LOGIC ;
		read		: IN STD_LOGIC ;
		reset		: IN STD_LOGIC ;
		busy		: OUT STD_LOGIC ;
		data_valid		: OUT STD_LOGIC ;
		dataout		: OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
		read_address		: OUT STD_LOGIC_VECTOR (23 DOWNTO 0)
	);
END asmicont;


ARCHITECTURE RTL OF asmicont IS

	ATTRIBUTE synthesis_clearbox: natural;
	ATTRIBUTE synthesis_clearbox OF RTL: ARCHITECTURE IS 2;
	ATTRIBUTE clearbox_macroname: string;
	ATTRIBUTE clearbox_macroname OF RTL: ARCHITECTURE IS "ALTASMI_PARALLEL";
	ATTRIBUTE clearbox_defparam: string;
	ATTRIBUTE clearbox_defparam OF RTL: ARCHITECTURE IS "data_width=STANDARD;epcs_type=EPCS64;intended_device_family=Cyclone V;lpm_hint=UNUSED;lpm_type=altasmi_parallel;page_size=1;port_bulk_erase=PORT_UNUSED;port_die_erase=PORT_UNUSED;port_en4b_addr=PORT_UNUSED;port_ex4b_addr=PORT_UNUSED;port_fast_read=PORT_UNUSED;port_illegal_erase=PORT_UNUSED;port_illegal_write=PORT_UNUSED;port_rdid_out=PORT_UNUSED;port_read_address=PORT_USED;port_read_dummyclk=PORT_UNUSED;port_read_rdid=PORT_UNUSED;port_read_sid=PORT_UNUSED;port_read_status=PORT_UNUSED;port_sector_erase=PORT_UNUSED;port_sector_protect=PORT_UNUSED;port_shift_bytes=PORT_UNUSED;port_wren=PORT_UNUSED;port_write=PORT_UNUSED;use_asmiblock=ON;use_eab=ON;write_dummy_clk=0;";
	SIGNAL sub_wire0	: STD_LOGIC ;
	SIGNAL sub_wire1	: STD_LOGIC ;
	SIGNAL sub_wire2	: STD_LOGIC_VECTOR (23 DOWNTO 0);
	SIGNAL sub_wire3	: STD_LOGIC_VECTOR (7 DOWNTO 0);



	COMPONENT asmicont_altasmi_parallel_qth2
	PORT (
			read	: IN STD_LOGIC ;
			addr	: IN STD_LOGIC_VECTOR (23 DOWNTO 0);
			busy	: OUT STD_LOGIC ;
			clkin	: IN STD_LOGIC ;
			data_valid	: OUT STD_LOGIC ;
			rden	: IN STD_LOGIC ;
			read_address	: OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
			reset	: IN STD_LOGIC ;
			dataout	: OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	busy    <= sub_wire0;
	data_valid    <= sub_wire1;
	read_address    <= sub_wire2(23 DOWNTO 0);
	dataout    <= sub_wire3(7 DOWNTO 0);

	asmicont_altasmi_parallel_qth2_component : asmicont_altasmi_parallel_qth2
	PORT MAP (
		read => read,
		addr => addr,
		clkin => clkin,
		rden => rden,
		reset => reset,
		busy => sub_wire0,
		data_valid => sub_wire1,
		read_address => sub_wire2,
		dataout => sub_wire3
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
-- Retrieval info: CONSTANT: DATA_WIDTH STRING "STANDARD"
-- Retrieval info: CONSTANT: EPCS_TYPE STRING "EPCS64"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
-- Retrieval info: CONSTANT: LPM_HINT STRING "UNUSED"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "altasmi_parallel"
-- Retrieval info: CONSTANT: PAGE_SIZE NUMERIC "1"
-- Retrieval info: CONSTANT: PORT_BULK_ERASE STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_DIE_ERASE STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_EN4B_ADDR STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_EX4B_ADDR STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_FAST_READ STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_ILLEGAL_ERASE STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_ILLEGAL_WRITE STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_RDID_OUT STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_READ_ADDRESS STRING "PORT_USED"
-- Retrieval info: CONSTANT: PORT_READ_DUMMYCLK STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_READ_RDID STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_READ_SID STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_READ_STATUS STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_SECTOR_ERASE STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_SECTOR_PROTECT STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_SHIFT_BYTES STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_WREN STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_WRITE STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: USE_ASMIBLOCK STRING "ON"
-- Retrieval info: CONSTANT: USE_EAB STRING "ON"
-- Retrieval info: CONSTANT: WRITE_DUMMY_CLK NUMERIC "0"
-- Retrieval info: USED_PORT: addr 0 0 24 0 INPUT NODEFVAL "addr[23..0]"
-- Retrieval info: CONNECT: @addr 0 0 24 0 addr 0 0 24 0
-- Retrieval info: USED_PORT: busy 0 0 0 0 OUTPUT NODEFVAL "busy"
-- Retrieval info: CONNECT: busy 0 0 0 0 @busy 0 0 0 0
-- Retrieval info: USED_PORT: clkin 0 0 0 0 INPUT NODEFVAL "clkin"
-- Retrieval info: CONNECT: @clkin 0 0 0 0 clkin 0 0 0 0
-- Retrieval info: USED_PORT: data_valid 0 0 0 0 OUTPUT NODEFVAL "data_valid"
-- Retrieval info: CONNECT: data_valid 0 0 0 0 @data_valid 0 0 0 0
-- Retrieval info: USED_PORT: dataout 0 0 8 0 OUTPUT NODEFVAL "dataout[7..0]"
-- Retrieval info: CONNECT: dataout 0 0 8 0 @dataout 0 0 8 0
-- Retrieval info: USED_PORT: rden 0 0 0 0 INPUT NODEFVAL "rden"
-- Retrieval info: CONNECT: @rden 0 0 0 0 rden 0 0 0 0
-- Retrieval info: USED_PORT: read 0 0 0 0 INPUT NODEFVAL "read"
-- Retrieval info: CONNECT: @read 0 0 0 0 read 0 0 0 0
-- Retrieval info: USED_PORT: read_address 0 0 24 0 OUTPUT NODEFVAL "read_address[23..0]"
-- Retrieval info: CONNECT: read_address 0 0 24 0 @read_address 0 0 24 0
-- Retrieval info: USED_PORT: reset 0 0 0 0 INPUT NODEFVAL "reset"
-- Retrieval info: CONNECT: @reset 0 0 0 0 reset 0 0 0 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL asmicont.vhd TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL asmicont.qip TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL asmicont.bsf TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL asmicont_inst.vhd TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL asmicont.inc TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL asmicont.cmp TRUE TRUE
